module up_memory(
	input	clk,
	input	nRst
);

endmodule
