module up_controller(
	input	clk,
	input	nRst
);

endmodule
