module up_reg_block(
	input	clk,
	input	nRst
);

endmodule
