module adc(
	input	clk,
	input	nRst,
   input [31:0] read
);

endmodule
