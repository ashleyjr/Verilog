module adc_tb;

	parameter CLK_PERIOD = 20;

	reg clk;
	reg nRst;
	reg [31:0] read;

	adc adc(
		.clk	(clk),
		.nRst	(nRst),
		.read	(read)
	);

	initial begin
		while(1) begin
			#(CLK_PERIOD/2) clk = 0;
			#(CLK_PERIOD/2) clk = 1;
		end	end

	initial begin
		$dumpfile("adc.vcd");
		$dumpvars(0,adc_tb);
	end

	initial begin
					nRst = 1;
		#100		nRst = 0;
		#100		nRst = 1;
		#1		read = 32'd2168958127;
		#1		read = 32'd2190430458;
		#1		read = 32'd2211898494;
		#1		read = 32'd2233360089;
		#1		read = 32'd2254813097;
		#1		read = 32'd2276255371;
		#1		read = 32'd2297684769;
		#1		read = 32'd2319099147;
		#1		read = 32'd2340496363;
		#1		read = 32'd2361874278;
		#1		read = 32'd2383230754;
		#1		read = 32'd2404563656;
		#1		read = 32'd2425870849;
		#1		read = 32'd2447150205;
		#1		read = 32'd2468399594;
		#1		read = 32'd2489616892;
		#1		read = 32'd2510799976;
		#1		read = 32'd2531946729;
		#1		read = 32'd2553055037;
		#1		read = 32'd2574122787;
		#1		read = 32'd2595147874;
		#1		read = 32'd2616128195;
		#1		read = 32'd2637061652;
		#1		read = 32'd2657946151;
		#1		read = 32'd2678779605;
		#1		read = 32'd2699559929;
		#1		read = 32'd2720285047;
		#1		read = 32'd2740952884;
		#1		read = 32'd2761561376;
		#1		read = 32'd2782108459;
		#1		read = 32'd2802592081;
		#1		read = 32'd2823010193;
		#1		read = 32'd2843360753;
		#1		read = 32'd2863641725;
		#1		read = 32'd2883851082;
		#1		read = 32'd2903986804;
		#1		read = 32'd2924046875;
		#1		read = 32'd2944029291;
		#1		read = 32'd2963932053;
		#1		read = 32'd2983753170;
		#1		read = 32'd3003490662;
		#1		read = 32'd3023142553;
		#1		read = 32'd3042706880;
		#1		read = 32'd3062181684;
		#1		read = 32'd3081565020;
		#1		read = 32'd3100854948;
		#1		read = 32'd3120049540;
		#1		read = 32'd3139146876;
		#1		read = 32'd3158145047;
		#1		read = 32'd3177042153;
		#1		read = 32'd3195836303;
		#1		read = 32'd3214525619;
		#1		read = 32'd3233108232;
		#1		read = 32'd3251582283;
		#1		read = 32'd3269945925;
		#1		read = 32'd3288197322;
		#1		read = 32'd3306334649;
		#1		read = 32'd3324356091;
		#1		read = 32'd3342259847;
		#1		read = 32'd3360044127;
		#1		read = 32'd3377707151;
		#1		read = 32'd3395247154;
		#1		read = 32'd3412662382;
		#1		read = 32'd3429951093;
		#1		read = 32'd3447111558;
		#1		read = 32'd3464142062;
		#1		read = 32'd3481040901;
		#1		read = 32'd3497806385;
		#1		read = 32'd3514436838;
		#1		read = 32'd3530930597;
		#1		read = 32'd3547286012;
		#1		read = 32'd3563501449;
		#1		read = 32'd3579575285;
		#1		read = 32'd3595505912;
		#1		read = 32'd3611291739;
		#1		read = 32'd3626931186;
		#1		read = 32'd3642422690;
		#1		read = 32'd3657764701;
		#1		read = 32'd3672955685;
		#1		read = 32'd3687994123;
		#1		read = 32'd3702878511;
		#1		read = 32'd3717607362;
		#1		read = 32'd3732179201;
		#1		read = 32'd3746592572;
		#1		read = 32'd3760846033;
		#1		read = 32'd3774938160;
		#1		read = 32'd3788867542;
		#1		read = 32'd3802632787;
		#1		read = 32'd3816232519;
		#1		read = 32'd3829665377;
		#1		read = 32'd3842930019;
		#1		read = 32'd3856025117;
		#1		read = 32'd3868949363;
		#1		read = 32'd3881701463;
		#1		read = 32'd3894280144;
		#1		read = 32'd3906684146;
		#1		read = 32'd3918912229;
		#1		read = 32'd3930963171;
		#1		read = 32'd3942835766;
		#1		read = 32'd3954528828;
		#1		read = 32'd3966041187;
		#1		read = 32'd3977371691;
		#1		read = 32'd3988519209;
		#1		read = 32'd3999482624;
		#1		read = 32'd4010260841;
		#1		read = 32'd4020852782;
		#1		read = 32'd4031257387;
		#1		read = 32'd4041473617;
		#1		read = 32'd4051500449;
		#1		read = 32'd4061336881;
		#1		read = 32'd4070981929;
		#1		read = 32'd4080434629;
		#1		read = 32'd4089694036;
		#1		read = 32'd4098759223;
		#1		read = 32'd4107629284;
		#1		read = 32'd4116303333;
		#1		read = 32'd4124780501;
		#1		read = 32'd4133059940;
		#1		read = 32'd4141140824;
		#1		read = 32'd4149022344;
		#1		read = 32'd4156703712;
		#1		read = 32'd4164184160;
		#1		read = 32'd4171462939;
		#1		read = 32'd4178539321;
		#1		read = 32'd4185412600;
		#1		read = 32'd4192082088;
		#1		read = 32'd4198547118;
		#1		read = 32'd4204807042;
		#1		read = 32'd4210861237;
		#1		read = 32'd4216709095;
		#1		read = 32'd4222350033;
		#1		read = 32'd4227783485;
		#1		read = 32'd4233008909;
		#1		read = 32'd4238025783;
		#1		read = 32'd4242833604;
		#1		read = 32'd4247431892;
		#1		read = 32'd4251820186;
		#1		read = 32'd4255998049;
		#1		read = 32'd4259965062;
		#1		read = 32'd4263720829;
		#1		read = 32'd4267264974;
		#1		read = 32'd4270597142;
		#1		read = 32'd4273717001;
		#1		read = 32'd4276624238;
		#1		read = 32'd4279318563;
		#1		read = 32'd4281799707;
		#1		read = 32'd4284067420;
		#1		read = 32'd4286121477;
		#1		read = 32'd4287961672;
		#1		read = 32'd4289587821;
		#1		read = 32'd4290999761;
		#1		read = 32'd4292197351;
		#1		read = 32'd4293180472;
		#1		read = 32'd4293949025;
		#1		read = 32'd4294502933;
		#1		read = 32'd4294842141;
		#1		read = 32'd4294966615;
		#1		read = 32'd4294876343;
		#1		read = 32'd4294571333;
		#1		read = 32'd4294051616;
		#1		read = 32'd4293317243;
		#1		read = 32'd4292368290;
		#1		read = 32'd4291204850;
		#1		read = 32'd4289827039;
		#1		read = 32'd4288234996;
		#1		read = 32'd4286428879;
		#1		read = 32'd4284408870;
		#1		read = 32'd4282175170;
		#1		read = 32'd4279728003;
		#1		read = 32'd4277067613;
		#1		read = 32'd4274194266;
		#1		read = 32'd4271108250;
		#1		read = 32'd4267809874;
		#1		read = 32'd4264299466;
		#1		read = 32'd4260577379;
		#1		read = 32'd4256643984;
		#1		read = 32'd4252499675;
		#1		read = 32'd4248144866;
		#1		read = 32'd4243579992;
		#1		read = 32'd4238805511;
		#1		read = 32'd4233821899;
		#1		read = 32'd4228629655;
		#1		read = 32'd4223229299;
		#1		read = 32'd4217621369;
		#1		read = 32'd4211806428;
		#1		read = 32'd4205785055;
		#1		read = 32'd4199557855;
		#1		read = 32'd4193125449;
		#1		read = 32'd4186488480;
		#1		read = 32'd4179647612;
		#1		read = 32'd4172603530;
		#1		read = 32'd4165356938;
		#1		read = 32'd4157908559;
		#1		read = 32'd4150259140;
		#1		read = 32'd4142409446;
		#1		read = 32'd4134360260;
		#1		read = 32'd4126112388;
		#1		read = 32'd4117666655;
		#1		read = 32'd4109023905;
		#1		read = 32'd4100185003;
		#1		read = 32'd4091150833;
		#1		read = 32'd4081922297;
		#1		read = 32'd4072500319;
		#1		read = 32'd4062885841;
		#1		read = 32'd4053079824;
		#1		read = 32'd4043083250;
		#1		read = 32'd4032897117;
		#1		read = 32'd4022522444;
		#1		read = 32'd4011960269;
		#1		read = 32'd4001211648;
		#1		read = 32'd3990277655;
		#1		read = 32'd3979159385;
		#1		read = 32'd3967857948;
		#1		read = 32'd3956374476;
		#1		read = 32'd3944710116;
		#1		read = 32'd3932866035;
		#1		read = 32'd3920843417;
		#1		read = 32'd3908643465;
		#1		read = 32'd3896267398;
		#1		read = 32'd3883716455;
		#1		read = 32'd3870991889;
		#1		read = 32'd3858094974;
		#1		read = 32'd3845027000;
		#1		read = 32'd3831789272;
		#1		read = 32'd3818383115;
		#1		read = 32'd3804809870;
		#1		read = 32'd3791070893;
		#1		read = 32'd3777167560;
		#1		read = 32'd3763101259;
		#1		read = 32'd3748873397;
		#1		read = 32'd3734485398;
		#1		read = 32'd3719938701;
		#1		read = 32'd3705234759;
		#1		read = 32'd3690375043;
		#1		read = 32'd3675361039;
		#1		read = 32'd3660194249;
		#1		read = 32'd3644876189;
		#1		read = 32'd3629408391;
		#1		read = 32'd3613792402;
		#1		read = 32'd3598029783;
		#1		read = 32'd3582122111;
		#1		read = 32'd3566070976;
		#1		read = 32'd3549877983;
		#1		read = 32'd3533544753;
		#1		read = 32'd3517072917;
		#1		read = 32'd3500464124;
		#1		read = 32'd3483720033;
		#1		read = 32'd3466842320;
		#1		read = 32'd3449832673;
		#1		read = 32'd3432692791;
		#1		read = 32'd3415424390;
		#1		read = 32'd3398029196;
		#1		read = 32'd3380508948;
		#1		read = 32'd3362865398;
		#1		read = 32'd3345100312;
		#1		read = 32'd3327215465;
		#1		read = 32'd3309212645;
		#1		read = 32'd3291093654;
		#1		read = 32'd3272860303;
		#1		read = 32'd3254514415;
		#1		read = 32'd3236057824;
		#1		read = 32'd3217492378;
		#1		read = 32'd3198819931;
		#1		read = 32'd3180042351;
		#1		read = 32'd3161161517;
		#1		read = 32'd3142179315;
		#1		read = 32'd3123097645;
		#1		read = 32'd3103918414;
		#1		read = 32'd3084643541;
		#1		read = 32'd3065274952;
		#1		read = 32'd3045814585;
		#1		read = 32'd3026264386;
		#1		read = 32'd3006626309;
		#1		read = 32'd2986902319;
		#1		read = 32'd2967094388;
		#1		read = 32'd2947204496;
		#1		read = 32'd2927234632;
		#1		read = 32'd2907186795;
		#1		read = 32'd2887062987;
		#1		read = 32'd2866865223;
		#1		read = 32'd2846595520;
		#1		read = 32'd2826255908;
		#1		read = 32'd2805848418;
		#1		read = 32'd2785375093;
		#1		read = 32'd2764837979;
		#1		read = 32'd2744239130;
		#1		read = 32'd2723580606;
		#1		read = 32'd2702864472;
		#1		read = 32'd2682092802;
		#1		read = 32'd2661267670;
		#1		read = 32'd2640391161;
		#1		read = 32'd2619465361;
		#1		read = 32'd2598492364;
		#1		read = 32'd2577474266;
		#1		read = 32'd2556413169;
		#1		read = 32'd2535311180;
		#1		read = 32'd2514170409;
		#1		read = 32'd2492992969;
		#1		read = 32'd2471780978;
		#1		read = 32'd2450536558;
		#1		read = 32'd2429261833;
		#1		read = 32'd2407958930;
		#1		read = 32'd2386629980;
		#1		read = 32'd2365277115;
		#1		read = 32'd2343902472;
		#1		read = 32'd2322508186;
		#1		read = 32'd2301096398;
		#1		read = 32'd2279669250;
		#1		read = 32'd2258228882;
		#1		read = 32'd2236777441;
		#1		read = 32'd2215317070;
		#1		read = 32'd2193849915;
		#1		read = 32'd2172378124;
		#1		read = 32'd2150903844;
		#1		read = 32'd2129429222;
		#1		read = 32'd2107956405;
		#1		read = 32'd2086487541;
		#1		read = 32'd2065024776;
		#1		read = 32'd2043570257;
		#1		read = 32'd2022126130;
		#1		read = 32'd2000694538;
		#1		read = 32'd1979277624;
		#1		read = 32'd1957877532;
		#1		read = 32'd1936496399;
		#1		read = 32'd1915136366;
		#1		read = 32'd1893799567;
		#1		read = 32'd1872488136;
		#1		read = 32'd1851204204;
		#1		read = 32'd1829949900;
		#1		read = 32'd1808727349;
		#1		read = 32'd1787538674;
		#1		read = 32'd1766385993;
		#1		read = 32'd1745271421;
		#1		read = 32'd1724197070;
		#1		read = 32'd1703165047;
		#1		read = 32'd1682177456;
		#1		read = 32'd1661236395;
		#1		read = 32'd1640343958;
		#1		read = 32'd1619502235;
		#1		read = 32'd1598713310;
		#1		read = 32'd1577979261;
		#1		read = 32'd1557302162;
		#1		read = 32'd1536684081;
		#1		read = 32'd1516127080;
		#1		read = 32'd1495633213;
		#1		read = 32'd1475204531;
		#1		read = 32'd1454843076;
		#1		read = 32'd1434550885;
		#1		read = 32'd1414329986;
		#1		read = 32'd1394182403;
		#1		read = 32'd1374110148;
		#1		read = 32'd1354115231;
		#1		read = 32'd1334199649;
		#1		read = 32'd1314365395;
		#1		read = 32'd1294614453;
		#1		read = 32'd1274948797;
		#1		read = 32'd1255370393;
		#1		read = 32'd1235881200;
		#1		read = 32'd1216483166;
		#1		read = 32'd1197178232;
		#1		read = 32'd1177968328;
		#1		read = 32'd1158855374;
		#1		read = 32'd1139841282;
		#1		read = 32'd1120927954;
		#1		read = 32'd1102117280;
		#1		read = 32'd1083411142;
		#1		read = 32'd1064811410;
		#1		read = 32'd1046319945;
		#1		read = 32'd1027938595;
		#1		read = 32'd1009669199;
		#1		read = 32'd991513584;
		#1		read = 32'd973473564;
		#1		read = 32'd955550944;
		#1		read = 32'd937747517;
		#1		read = 32'd920065062;
		#1		read = 32'd902505348;
		#1		read = 32'd885070131;
		#1		read = 32'd867761154;
		#1		read = 32'd850580149;
		#1		read = 32'd833528832;
		#1		read = 32'd816608910;
		#1		read = 32'd799822075;
		#1		read = 32'd783170004;
		#1		read = 32'd766654364;
		#1		read = 32'd750276805;
		#1		read = 32'd734038966;
		#1		read = 32'd717942470;
		#1		read = 32'd701988928;
		#1		read = 32'd686179933;
		#1		read = 32'd670517068;
		#1		read = 32'd655001898;
		#1		read = 32'd639635974;
		#1		read = 32'd624420835;
		#1		read = 32'd609358000;
		#1		read = 32'd594448977;
		#1		read = 32'd579695256;
		#1		read = 32'd565098312;
		#1		read = 32'd550659606;
		#1		read = 32'd536380581;
		#1		read = 32'd522262665;
		#1		read = 32'd508307269;
		#1		read = 32'd494515790;
		#1		read = 32'd480889606;
		#1		read = 32'd467430080;
		#1		read = 32'd454138558;
		#1		read = 32'd441016369;
		#1		read = 32'd428064826;
		#1		read = 32'd415285223;
		#1		read = 32'd402678838;
		#1		read = 32'd390246932;
		#1		read = 32'd377990749;
		#1		read = 32'd365911513;
		#1		read = 32'd354010434;
		#1		read = 32'd342288700;
		#1		read = 32'd330747483;
		#1		read = 32'd319387940;
		#1		read = 32'd308211204;
		#1		read = 32'd297218393;
		#1		read = 32'd286410608;
		#1		read = 32'd275788929;
		#1		read = 32'd265354417;
		#1		read = 32'd255108117;
		#1		read = 32'd245051053;
		#1		read = 32'd235184230;
		#1		read = 32'd225508636;
		#1		read = 32'd216025238;
		#1		read = 32'd206734984;
		#1		read = 32'd197638803;
		#1		read = 32'd188737605;
		#1		read = 32'd180032280;
		#1		read = 32'd171523698;
		#1		read = 32'd163212711;
		#1		read = 32'd155100150;
		#1		read = 32'd147186825;
		#1		read = 32'd139473528;
		#1		read = 32'd131961030;
		#1		read = 32'd124650083;
		#1		read = 32'd117541418;
		#1		read = 32'd110635745;
		#1		read = 32'd103933755;
		#1		read = 32'd97436118;
		#1		read = 32'd91143485;
		#1		read = 32'd85056484;
		#1		read = 32'd79175724;
		#1		read = 32'd73501793;
		#1		read = 32'd68035258;
		#1		read = 32'd62776667;
		#1		read = 32'd57726544;
		#1		read = 32'd52885395;
		#1		read = 32'd48253705;
		#1		read = 32'd43831936;
		#1		read = 32'd39620530;
		#1		read = 32'd35619909;
		#1		read = 32'd31830472;
		#1		read = 32'd28252599;
		#1		read = 32'd24886647;
		#1		read = 32'd21732953;
		#1		read = 32'd18791833;
		#1		read = 32'd16063579;
		#1		read = 32'd13548467;
		#1		read = 32'd11246745;
		#1		read = 32'd9158646;
		#1		read = 32'd7284378;
		#1		read = 32'd5624127;
		#1		read = 32'd4178061;
		#1		read = 32'd2946323;
		#1		read = 32'd1929038;
		#1		read = 32'd1126306;
		#1		read = 32'd538208;
		#1		read = 32'd164803;
		#1		read = 32'd6128;
		#1		read = 32'd62199;
		#1		read = 32'd333010;
		#1		read = 32'd818535;
		#1		read = 32'd1518724;
		#1		read = 32'd2433508;
		#1		read = 32'd3562795;
		#1		read = 32'd4906473;
		#1		read = 32'd6464406;
		#1		read = 32'd8236440;
		#1		read = 32'd10222396;
		#1		read = 32'd12422077;
		#1		read = 32'd14835262;
		#1		read = 32'd17461711;
		#1		read = 32'd20301159;
		#1		read = 32'd23353325;
		#1		read = 32'd26617901;
		#1		read = 32'd30094562;
		#1		read = 32'd33782961;
		#1		read = 32'd37682727;
		#1		read = 32'd41793473;
		#1		read = 32'd46114785;
		#1		read = 32'd50646232;
		#1		read = 32'd55387362;
		#1		read = 32'd60337699;
		#1		read = 32'd65496749;
		#1		read = 32'd70863996;
		#1		read = 32'd76438904;
		#1		read = 32'd82220914;
		#1		read = 32'd88209448;
		#1		read = 32'd94403909;
		#1		read = 32'd100803676;
		#1		read = 32'd107408108;
		#1		read = 32'd114216547;
		#1		read = 32'd121228311;
		#1		read = 32'd128442699;
		#1		read = 32'd135858989;
		#1		read = 32'd143476440;
		#1		read = 32'd151294289;
		#1		read = 32'd159311757;
		#1		read = 32'd167528039;
		#1		read = 32'd175942316;
		#1		read = 32'd184553745;
		#1		read = 32'd193361465;
		#1		read = 32'd202364597;
		#1		read = 32'd211562238;
		#1		read = 32'd220953470;
		#1		read = 32'd230537353;
		#1		read = 32'd240312929;
		#1		read = 32'd250279221;
		#1		read = 32'd260435232;
		#1		read = 32'd270779946;
		#1		read = 32'd281312328;
		#1		read = 32'd292031327;
		#1		read = 32'd302935869;
		#1		read = 32'd314024864;
		#1		read = 32'd325297203;
		#1		read = 32'd336751760;
		#1		read = 32'd348387389;
		#1		read = 32'd360202925;
		#1		read = 32'd372197188;
		#1		read = 32'd384368978;
		#1		read = 32'd396717079;
		#1		read = 32'd409240254;
		#1		read = 32'd421937252;
		#1		read = 32'd434806804;
		#1		read = 32'd447847622;
		#1		read = 32'd461058402;
		#1		read = 32'd474437823;
		#1		read = 32'd487984547;
		#1		read = 32'd501697220;
		#1		read = 32'd515574470;
		#1		read = 32'd529614910;
		#1		read = 32'd543817135;
		#1		read = 32'd558179725;
		#1		read = 32'd572701245;
		#1		read = 32'd587380242;
		#1		read = 32'd602215247;
		#1		read = 32'd617204778;
		#1		read = 32'd632347336;
		#1		read = 32'd647641406;
		#1		read = 32'd663085459;
		#1		read = 32'd678677951;
		#1		read = 32'd694417322;
		#1		read = 32'd710301998;
		#1		read = 32'd726330391;
		#1		read = 32'd742500899;
		#1		read = 32'd758811903;
		#1		read = 32'd775261774;
		#1		read = 32'd791848866;
		#1		read = 32'd808571520;
		#1		read = 32'd825428064;
		#1		read = 32'd842416812;
		#1		read = 32'd859536066;
		#1		read = 32'd876784114;
		#1		read = 32'd894159231;
		#1		read = 32'd911659679;
		#1		read = 32'd929283709;
		#1		read = 32'd947029557;
		#1		read = 32'd964895450;
		#1		read = 32'd982879601;
		#1		read = 32'd1000980211;
		#1		read = 32'd1019195471;
		#1		read = 32'd1037523558;
		#1		read = 32'd1055962640;
		#1		read = 32'd1074510874;
		#1		read = 32'd1093166404;
		#1		read = 32'd1111927365;
		#1		read = 32'd1130791881;
		#1		read = 32'd1149758065;
		#1		read = 32'd1168824021;
		#1		read = 32'd1187987842;
		#1		read = 32'd1207247611;
		#1		read = 32'd1226601404;
		#1		read = 32'd1246047284;
		#1		read = 32'd1265583307;
		#1		read = 32'd1285207519;
		#1		read = 32'd1304917958;
		#1		read = 32'd1324712653;
		#1		read = 32'd1344589624;
		#1		read = 32'd1364546884;
		#1		read = 32'd1384582437;
		#1		read = 32'd1404694280;
		#1		read = 32'd1424880400;
		#1		read = 32'd1445138781;
		#1		read = 32'd1465467396;
		#1		read = 32'd1485864211;
		#1		read = 32'd1506327188;
		#1		read = 32'd1526854280;
		#1		read = 32'd1547443435;
		#1		read = 32'd1568092593;
		#1		read = 32'd1588799689;
		#1		read = 32'd1609562654;
		#1		read = 32'd1630379410;
		#1		read = 32'd1651247876;
		#1		read = 32'd1672165966;
		#1		read = 32'd1693131586;
		#1		read = 32'd1714142642;
		#1		read = 32'd1735197031;
		#1		read = 32'd1756292649;
		#1		read = 32'd1777427385;
		#1		read = 32'd1798599127;
		#1		read = 32'd1819805757;
		#1		read = 32'd1841045154;
		#1		read = 32'd1862315195;
		#1		read = 32'd1883613753;
		#1		read = 32'd1904938697;
		#1		read = 32'd1926287896;
		#1		read = 32'd1947659214;
		#1		read = 32'd1969050514;
		#1		read = 32'd1990459658;
		#1		read = 32'd2011884503;
		#1		read = 32'd2033322909;
		#1		read = 32'd2054772730;
		#1		read = 32'd2076231823;
		#1		read = 32'd2097698041;
		#1		read = 32'd2119169237;
		#1		read = 32'd2140643264;
		#1		read = 32'd2162117976;
		#1		read = 32'd2183591224;
		#1		read = 32'd2205060862;
		#1		read = 32'd2226524742;
		#1		read = 32'd2247980717;
		#1		read = 32'd2269426644;
		#1		read = 32'd2290860376;
		#1		read = 32'd2312279770;
		#1		read = 32'd2333682685;
		#1		read = 32'd2355066980;
		#1		read = 32'd2376430517;
		#1		read = 32'd2397771160;
		#1		read = 32'd2419086774;
		#1		read = 32'd2440375227;
		#1		read = 32'd2461634392;
		#1		read = 32'd2482862143;
		#1		read = 32'd2504056355;
		#1		read = 32'd2525214911;
		#1		read = 32'd2546335694;
		#1		read = 32'd2567416592;
		#1		read = 32'd2588455497;
		#1		read = 32'd2609450305;
		#1		read = 32'd2630398917;
		#1		read = 32'd2651299237;
		#1		read = 32'd2672149177;
		#1		read = 32'd2692946651;
		#1		read = 32'd2713689578;
		#1		read = 32'd2734375886;
		#1		read = 32'd2755003505;
		#1		read = 32'd2775570372;
		#1		read = 32'd2796074431;
		#1		read = 32'd2816513632;
		#1		read = 32'd2836885930;
		#1		read = 32'd2857189289;
		#1		read = 32'd2877421677;
		#1		read = 32'd2897581073;
		#1		read = 32'd2917665459;
		#1		read = 32'd2937672828;
		#1		read = 32'd2957601178;
		#1		read = 32'd2977448517;
		#1		read = 32'd2997212861;
		#1		read = 32'd3016892232;
		#1		read = 32'd3036484664;
		#1		read = 32'd3055988196;
		#1		read = 32'd3075400878;
		#1		read = 32'd3094720769;
		#1		read = 32'd3113945937;
		#1		read = 32'd3133074460;
		#1		read = 32'd3152104425;
		#1		read = 32'd3171033928;
		#1		read = 32'd3189861077;
		#1		read = 32'd3208583990;
		#1		read = 32'd3227200793;
		#1		read = 32'd3245709625;
		#1		read = 32'd3264108636;
		#1		read = 32'd3282395985;
		#1		read = 32'd3300569844;
		#1		read = 32'd3318628395;
		#1		read = 32'd3336569833;
		#1		read = 32'd3354392363;
		#1		read = 32'd3372094203;
		#1		read = 32'd3389673583;
		#1		read = 32'd3407128746;
		#1		read = 32'd3424457944;
		#1		read = 32'd3441659447;
		#1		read = 32'd3458731533;
		#1		read = 32'd3475672495;
		#1		read = 32'd3492480639;
		#1		read = 32'd3509154285;
		#1		read = 32'd3525691765;
		#1		read = 32'd3542091425;
		#1		read = 32'd3558351626;
		#1		read = 32'd3574470741;
		#1		read = 32'd3590447158;
		#1		read = 32'd3606279280;
		#1		read = 32'd3621965524;
		#1		read = 32'd3637504321;
		#1		read = 32'd3652894118;
		#1		read = 32'd3668133374;
		#1		read = 32'd3683220567;
		#1		read = 32'd3698154187;
		#1		read = 32'd3712932742;
		#1		read = 32'd3727554752;
		#1		read = 32'd3742018758;
		#1		read = 32'd3756323311;
		#1		read = 32'd3770466981;
		#1		read = 32'd3784448354;
		#1		read = 32'd3798266032;
		#1		read = 32'd3811918634;
		#1		read = 32'd3825404793;
		#1		read = 32'd3838723162;
		#1		read = 32'd3851872408;
		#1		read = 32'd3864851216;
		#1		read = 32'd3877658289;
		#1		read = 32'd3890292346;
		#1		read = 32'd3902752124;
		#1		read = 32'd3915036377;
		#1		read = 32'd3927143875;
		#1		read = 32'd3939073409;
		#1		read = 32'd3950823786;
		#1		read = 32'd3962393830;
		#1		read = 32'd3973782384;
		#1		read = 32'd3984988311;
		#1		read = 32'd3996010488;
		#1		read = 32'd4006847814;
		#1		read = 32'd4017499205;
		#1		read = 32'd4027963597;
		#1		read = 32'd4038239941;
		#1		read = 32'd4048327212;
		#1		read = 32'd4058224400;
		#1		read = 32'd4067930516;
		#1		read = 32'd4077444588;
		#1		read = 32'd4086765666;
		#1		read = 32'd4095892817;
		#1		read = 32'd4104825129;
		#1		read = 32'd4113561709;
		#1		read = 32'd4122101682;
		#1		read = 32'd4130444196;
		#1		read = 32'd4138588414;
		#1		read = 32'd4146533524;
		#1		read = 32'd4154278731;
		#1		read = 32'd4161823260;
		#1		read = 32'd4169166357;
		#1		read = 32'd4176307286;
		#1		read = 32'd4183245336;
		#1		read = 32'd4189979811;
		#1		read = 32'd4196510038;
		#1		read = 32'd4202835364;
		#1		read = 32'd4208955156;
		#1		read = 32'd4214868803;
		#1		read = 32'd4220575713;
		#1		read = 32'd4226075316;
		#1		read = 32'd4231367062;
		#1		read = 32'd4236450420;
		#1		read = 32'd4241324884;
		#1		read = 32'd4245989966;
		#1		read = 32'd4250445198;
		#1		read = 32'd4254690137;
		#1		read = 32'd4258724356;
		#1		read = 32'd4262547453;
		#1		read = 32'd4266159045;
		#1		read = 32'd4269558772;
		#1		read = 32'd4272746293;
		#1		read = 32'd4275721289;
		#1		read = 32'd4278483463;
		#1		read = 32'd4281032539;
		#1		read = 32'd4283368262;
		#1		read = 32'd4285490399;
		#1		read = 32'd4287398736;
		#1		read = 32'd4289093084;
		#1		read = 32'd4290573273;
		#1		read = 32'd4291839154;
		#1		read = 32'd4292890602;
		#1		read = 32'd4293727510;
		#1		read = 32'd4294349797;
		#1		read = 32'd4294757398;
		#1		read = 32'd4294950274;
		#1		read = 32'd4294928404;
		#1		read = 32'd4294691793;
		#1		read = 32'd4294240462;
		#1		read = 32'd4293574457;
		#1		read = 32'd4292693845;
		#1		read = 32'd4291598714;
		#1		read = 32'd4290289173;
		#1		read = 32'd4288765353;
		#1		read = 32'd4287027407;
		#1		read = 32'd4285075508;
		#1		read = 32'd4282909852;
		#1		read = 32'd4280530655;
		#1		read = 32'd4277938155;
		#1		read = 32'd4275132611;
		#1		read = 32'd4272114305;
		#1		read = 32'd4268883537;
		#1		read = 32'd4265440630;
		#1		read = 32'd4261785930;
		#1		read = 32'd4257919802;
		#1		read = 32'd4253842631;
		#1		read = 32'd4249554827;
		#1		read = 32'd4245056817;
		#1		read = 32'd4240349051;
		#1		read = 32'd4235432001;
		#1		read = 32'd4230306157;
		#1		read = 32'd4224972033;
		#1		read = 32'd4219430162;
		#1		read = 32'd4213681098;
		#1		read = 32'd4207725416;
		#1		read = 32'd4201563712;
		#1		read = 32'd4195196601;
		#1		read = 32'd4188624720;
		#1		read = 32'd4181848728;
		#1		read = 32'd4174869300;
		#1		read = 32'd4167687136;
		#1		read = 32'd4160302953;
		#1		read = 32'd4152717489;
		#1		read = 32'd4144931504;
		#1		read = 32'd4136945776;
		#1		read = 32'd4128761103;
		#1		read = 32'd4120378304;
		#1		read = 32'd4111798218;
		#1		read = 32'd4103021701;
		#1		read = 32'd4094049632;
		#1		read = 32'd4084882909;
		#1		read = 32'd4075522447;
		#1		read = 32'd4065969182;
		#1		read = 32'd4056224071;
		#1		read = 32'd4046288088;
		#1		read = 32'd4036162225;
		#1		read = 32'd4025847496;
		#1		read = 32'd4015344933;
		#1		read = 32'd4004655585;
		#1		read = 32'd3993780521;
		#1		read = 32'd3982720829;
		#1		read = 32'd3971477615;
		#1		read = 32'd3960052003;
		#1		read = 32'd3948445135;
		#1		read = 32'd3936658173;
		#1		read = 32'd3924692295;
		#1		read = 32'd3912548698;
		#1		read = 32'd3900228595;
		#1		read = 32'd3887733220;
		#1		read = 32'd3875063821;
		#1		read = 32'd3862221665;
		#1		read = 32'd3849208038;
		#1		read = 32'd3836024239;
		#1		read = 32'd3822671587;
		#1		read = 32'd3809151418;
		#1		read = 32'd3795465084;
		#1		read = 32'd3781613953;
		#1		read = 32'd3767599410;
		#1		read = 32'd3753422857;
		#1		read = 32'd3739085711;
		#1		read = 32'd3724589407;
		#1		read = 32'd3709935393;
		#1		read = 32'd3695125135;
		#1		read = 32'd3680160115;
		#1		read = 32'd3665041828;
		#1		read = 32'd3649771787;
		#1		read = 32'd3634351518;
		#1		read = 32'd3618782563;
		#1		read = 32'd3603066480;
		#1		read = 32'd3587204840;
		#1		read = 32'd3571199229;
		#1		read = 32'd3555051247;
		#1		read = 32'd3538762510;
		#1		read = 32'd3522334646;
		#1		read = 32'd3505769298;
		#1		read = 32'd3489068123;
		#1		read = 32'd3472232791;
		#1		read = 32'd3455264984;
		#1		read = 32'd3438166401;
		#1		read = 32'd3420938750;
		#1		read = 32'd3403583755;
		#1		read = 32'd3386103151;
		#1		read = 32'd3368498686;
		#1		read = 32'd3350772121;
		#1		read = 32'd3332925227;
		#1		read = 32'd3314959791;
		#1		read = 32'd3296877608;
		#1		read = 32'd3278680486;
		#1		read = 32'd3260370246;
		#1		read = 32'd3241948718;
		#1		read = 32'd3223417745;
		#1		read = 32'd3204779178;
		#1		read = 32'd3186034884;
		#1		read = 32'd3167186735;
		#1		read = 32'd3148236616;
		#1		read = 32'd3129186423;
		#1		read = 32'd3110038061;
		#1		read = 32'd3090793444;
		#1		read = 32'd3071454496;
		#1		read = 32'd3052023153;
		#1		read = 32'd3032501356;
		#1		read = 32'd3012891058;
		#1		read = 32'd2993194220;
		#1		read = 32'd2973412812;
		#1		read = 32'd2953548812;
		#1		read = 32'd2933604206;
		#1		read = 32'd2913580988;
		#1		read = 32'd2893481161;
		#1		read = 32'd2873306735;
		#1		read = 32'd2853059728;
		#1		read = 32'd2832742163;
		#1		read = 32'd2812356073;
		#1		read = 32'd2791903497;
		#1		read = 32'd2771386479;
		#1		read = 32'd2750807071;
		#1		read = 32'd2730167331;
		#1		read = 32'd2709469324;
		#1		read = 32'd2688715118;
		#1		read = 32'd2667906790;
		#1		read = 32'd2647046420;
		#1		read = 32'd2626136094;
		#1		read = 32'd2605177903;
		#1		read = 32'd2584173943;
		#1		read = 32'd2563126314;
		#1		read = 32'd2542037122;
		#1		read = 32'd2520908474;
		#1		read = 32'd2499742485;
		#1		read = 32'd2478541269;
		#1		read = 32'd2457306949;
		#1		read = 32'd2436041646;
		#1		read = 32'd2414747487;
		#1		read = 32'd2393426603;
		#1		read = 32'd2372081124;
		#1		read = 32'd2350713186;
		#1		read = 32'd2329324925;
		#1		read = 32'd2307918480;
		#1		read = 32'd2286495992;
		#1		read = 32'd2265059602;
		#1		read = 32'd2243611455;
		#1		read = 32'd2222153696;
		#1		read = 32'd2200688469;
		#1		read = 32'd2179217922;
		#1		read = 32'd2157744202;
		#1		read = 32'd2136269455;
		#1		read = 32'd2114795830;
		#1		read = 32'd2093325474;
		#1		read = 32'd2071860533;
		#1		read = 32'd2050403155;
		#1		read = 32'd2028955485;
		#1		read = 32'd2007519667;
		#1		read = 32'd1986097846;
		#1		read = 32'd1964692163;
		#1		read = 32'd1943304759;
		#1		read = 32'd1921937773;
		#1		read = 32'd1900593341;
		#1		read = 32'd1879273598;
		#1		read = 32'd1857980676;
		#1		read = 32'd1836716704;
		#1		read = 32'd1815483808;
		#1		read = 32'd1794284112;
		#1		read = 32'd1773119736;
		#1		read = 32'd1751992796;
		#1		read = 32'd1730905404;
		#1		read = 32'd1709859670;
		#1		read = 32'd1688857698;
		#1		read = 32'd1667901589;
		#1		read = 32'd1646993437;
		#1		read = 32'd1626135333;
		#1		read = 32'd1605329364;
		#1		read = 32'd1584577610;
		#1		read = 32'd1563882147;
		#1		read = 32'd1543245042;
		#1		read = 32'd1522668362;
		#1		read = 32'd1502154162;
		#1		read = 32'd1481704494;
		#1		read = 32'd1461321404;
		#1		read = 32'd1441006930;
		#1		read = 32'd1420763103;
		#1		read = 32'd1400591947;
		#1		read = 32'd1380495480;
		#1		read = 32'd1360475711;
		#1		read = 32'd1340534642;
		#1		read = 32'd1320674267;
		#1		read = 32'd1300896572;
		#1		read = 32'd1281203536;
		#1		read = 32'd1261597127;
		#1		read = 32'd1242079305;
		#1		read = 32'd1222652024;
		#1		read = 32'd1203317225;
		#1		read = 32'd1184076841;
		#1		read = 32'd1164932798;
		#1		read = 32'd1145887009;
		#1		read = 32'd1126941378;
		#1		read = 32'd1108097801;
		#1		read = 32'd1089358162;
		#1		read = 32'd1070724334;
		#1		read = 32'd1052198182;
		#1		read = 32'd1033781557;
		#1		read = 32'd1015476301;
		#1		read = 32'd997284245;
		#1		read = 32'd979207208;
		#1		read = 32'd961246998;
		#1		read = 32'd943405410;
		#1		read = 32'd925684230;
		#1		read = 32'd908085228;
		#1		read = 32'd890610165;
		#1		read = 32'd873260788;
		#1		read = 32'd856038833;
		#1		read = 32'd838946021;
		#1		read = 32'd821984061;
		#1		read = 32'd805154651;
		#1		read = 32'd788459472;
		#1		read = 32'd771900194;
		#1		read = 32'd755478474;
		#1		read = 32'd739195953;
		#1		read = 32'd723054260;
		#1		read = 32'd707055008;
		#1		read = 32'd691199798;
		#1		read = 32'd675490216;
		#1		read = 32'd659927831;
		#1		read = 32'd644514201;
		#1		read = 32'd629250866;
		#1		read = 32'd614139354;
		#1		read = 32'd599181174;
		#1		read = 32'd584377824;
		#1		read = 32'd569730782;
		#1		read = 32'd555241515;
		#1		read = 32'd540911471;
		#1		read = 32'd526742082;
		#1		read = 32'd512734767;
		#1		read = 32'd498890925;
		#1		read = 32'd485211941;
		#1		read = 32'd471699182;
		#1		read = 32'd458354001;
		#1		read = 32'd445177731;
		#1		read = 32'd432171690;
		#1		read = 32'd419337179;
		#1		read = 32'd406675482;
		#1		read = 32'd394187863;
		#1		read = 32'd381875573;
		#1		read = 32'd369739842;
		#1		read = 32'd357781884;
		#1		read = 32'd346002895;
		#1		read = 32'd334404052;
		#1		read = 32'd322986516;
		#1		read = 32'd311751428;
		#1		read = 32'd300699912;
		#1		read = 32'd289833072;
		#1		read = 32'd279151996;
		#1		read = 32'd268657752;
		#1		read = 32'd258351388;
		#1		read = 32'd248233937;
		#1		read = 32'd238306408;
		#1		read = 32'd228569796;
		#1		read = 32'd219025073;
		#1		read = 32'd209673195;
		#1		read = 32'd200515097;
		#1		read = 32'd191551693;
		#1		read = 32'd182783881;
		#1		read = 32'd174212537;
		#1		read = 32'd165838519;
		#1		read = 32'd157662664;
		#1		read = 32'd149685789;
		#1		read = 32'd141908692;
		#1		read = 32'd134332152;
		#1		read = 32'd126956924;
		#1		read = 32'd119783748;
		#1		read = 32'd112813340;
		#1		read = 32'd106046397;
		#1		read = 32'd99483596;
		#1		read = 32'd93125593;
		#1		read = 32'd86973025;
		#1		read = 32'd81026506;
		#1		read = 32'd75286631;
		#1		read = 32'd69753974;
		#1		read = 32'd64429088;
		#1		read = 32'd59312506;
		#1		read = 32'd54404739;
		#1		read = 32'd49706279;
		#1		read = 32'd45217594;
		#1		read = 32'd40939134;
		#1		read = 32'd36871327;
		#1		read = 32'd33014580;
		#1		read = 32'd29369277;
		#1		read = 32'd25935784;
		#1		read = 32'd22714445;
		#1		read = 32'd19705580;
		#1		read = 32'd16909491;
		#1		read = 32'd14326458;
		#1		read = 32'd11956739;
		#1		read = 32'd9800571;
		#1		read = 32'd7858170;
		#1		read = 32'd6129729;
		#1		read = 32'd4615422;
		#1		read = 32'd3315400;
		#1		read = 32'd2229793;
		#1		read = 32'd1358709;
		#1		read = 32'd702236;
		#1		read = 32'd260440;
		#1		read = 32'd33364;
		#1		read = 32'd21031;
		#1		read = 32'd223443;
		#1		read = 32'd640579;
		#1		read = 32'd1272398;
		#1		read = 32'd2118836;
		#1		read = 32'd3179808;
		#1		read = 32'd4455209;
		#1		read = 32'd5944911;
		#1		read = 32'd7648766;
		#1		read = 32'd9566602;
		#1		read = 32'd11698228;
		#1		read = 32'd14043430;
		#1		read = 32'd16601975;
		#1		read = 32'd19373607;
		#1		read = 32'd22358047;
		#1		read = 32'd25554999;
		#1		read = 32'd28964141;
		#1		read = 32'd32585134;
		#1		read = 32'd36417615;
		#1		read = 32'd40461200;
		#1		read = 32'd44715486;
		#1		read = 32'd49180047;
		#1		read = 32'd53854437;
		#1		read = 32'd58738188;
		#1		read = 32'd63830812;
		#1		read = 32'd69131799;
		#1		read = 32'd74640620;
		#1		read = 32'd80356723;
		#1		read = 32'd86279537;
		#1		read = 32'd92408470;
		#1		read = 32'd98742909;
		#1		read = 32'd105282220;
		#1		read = 32'd112025750;
		#1		read = 32'd118972823;
		#1		read = 32'd126122746;
		#1		read = 32'd133474804;
		#1		read = 32'd141028261;
		#1		read = 32'd148782361;
		#1		read = 32'd156736330;
		#1		read = 32'd164889372;
		#1		read = 32'd173240672;
		#1		read = 32'd181789394;
		#1		read = 32'd190534685;
		#1		read = 32'd199475668;
		#1		read = 32'd208611451;
		#1		read = 32'd217941119;
		#1		read = 32'd227463740;
		#1		read = 32'd237178362;
		#1		read = 32'd247084012;
		#1		read = 32'd257179701;
		#1		read = 32'd267464418;
		#1		read = 32'd277937136;
		#1		read = 32'd288596807;
		#1		read = 32'd299442365;
		#1		read = 32'd310472726;
		#1		read = 32'd321686786;
		#1		read = 32'd333083424;
		#1		read = 32'd344661501;
		#1		read = 32'd356419859;
		#1		read = 32'd368357322;
		#1		read = 32'd380472695;
		#1		read = 32'd392764768;
		#1		read = 32'd405232312;
		#1		read = 32'd417874080;
		#1		read = 32'd430688806;
		#1		read = 32'd443675211;
		#1		read = 32'd456831996;
		#1		read = 32'd470157844;
		#1		read = 32'd483651423;
		#1		read = 32'd497311384;
		#1		read = 32'd511136361;
		#1		read = 32'd525124972;
		#1		read = 32'd539275817;
		#1		read = 32'd553587481;
		#1		read = 32'd568058534;
		#1		read = 32'd582687528;
		#1		read = 32'd597473000;
		#1		read = 32'd612413472;
		#1		read = 32'd627507449;
		#1		read = 32'd642753423;
		#1		read = 32'd658149869;
		#1		read = 32'd673695247;
		#1		read = 32'd689388002;
		#1		read = 32'd705226566;
		#1		read = 32'd721209355;
		#1		read = 32'd737334769;
		#1		read = 32'd753601198;
		#1		read = 32'd770007013;
		#1		read = 32'd786550575;
		#1		read = 32'd803230229;
		#1		read = 32'd820044307;
		#1		read = 32'd836991128;
		#1		read = 32'd854068998;
		#1		read = 32'd871276207;
		#1		read = 32'd888611037;
		#1		read = 32'd906071752;
		#1		read = 32'd923656608;
		#1		read = 32'd941363845;
		#1		read = 32'd959191694;
		#1		read = 32'd977138370;
		#1		read = 32'd995202081;
		#1		read = 32'd1013381018;
		#1		read = 32'd1031673365;
		#1		read = 32'd1050077291;
		#1		read = 32'd1068590958;
		#1		read = 32'd1087212513;
		#1		read = 32'd1105940094;
		#1		read = 32'd1124771828;
		#1		read = 32'd1143705833;
		#1		read = 32'd1162740215;
		#1		read = 32'd1181873071;
		#1		read = 32'd1201102486;
		#1		read = 32'd1220426539;
		#1		read = 32'd1239843297;
		#1		read = 32'd1259350818;
		#1		read = 32'd1278947152;
		#1		read = 32'd1298630339;
		#1		read = 32'd1318398410;
		#1		read = 32'd1338249389;
		#1		read = 32'd1358181291;
		#1		read = 32'd1378192122;
		#1		read = 32'd1398279882;
		#1		read = 32'd1418442562;
		#1		read = 32'd1438678145;
		#1		read = 32'd1458984608;
		#1		read = 32'd1479359921;
		#1		read = 32'd1499802045;
		#1		read = 32'd1520308937;
		#1		read = 32'd1540878546;
		#1		read = 32'd1561508815;
		#1		read = 32'd1582197680;
		#1		read = 32'd1602943074;
		#1		read = 32'd1623742922;
		#1		read = 32'd1644595143;
		#1		read = 32'd1665497653;
		#1		read = 32'd1686448361;
		#1		read = 32'd1707445172;
		#1		read = 32'd1728485986;
		#1		read = 32'd1749568700;
		#1		read = 32'd1770691205;
		#1		read = 32'd1791851389;
		#1		read = 32'd1813047136;
		#1		read = 32'd1834276326;
		#1		read = 32'd1855536837;
		#1		read = 32'd1876826542;
		#1		read = 32'd1898143313;
		#1		read = 32'd1919485018;
		#1		read = 32'd1940849522;
		#1		read = 32'd1962234689;
		#1		read = 32'd1983638381;
		#1		read = 32'd2005058458;
		#1		read = 32'd2026492777;
		#1		read = 32'd2047939195;
		#1		read = 32'd2069395567;
		#1		read = 32'd2090859748;
		#1		read = 32'd2112329592;
		#1		read = 32'd2133802950;
		#1		read = 32'd2155277677;
		#1		read = 32'd2176751625;
		#1		read = 32'd2198222645;
		#1		read = 32'd2219688592;
		#1		read = 32'd2241147318;
		#1		read = 32'd2262596679;
		#1		read = 32'd2284034527;
		#1		read = 32'd2305458721;
		#1		read = 32'd2326867118;
		#1		read = 32'd2348257576;
		#1		read = 32'd2369627957;
		#1		read = 32'd2390976124;
		#1		read = 32'd2412299942;
		#1		read = 32'd2433597278;
		#1		read = 32'd2454866004;
		#1		read = 32'd2476103991;
		#1		read = 32'd2497309116;
		#1		read = 32'd2518479260;
		#1		read = 32'd2539612304;
		#1		read = 32'd2560706135;
		#1		read = 32'd2581758645;
		#1		read = 32'd2602767727;
		#1		read = 32'd2623731282;
		#1		read = 32'd2644647212;
		#1		read = 32'd2665513426;
		#1		read = 32'd2686327837;
		#1		read = 32'd2707088365;
		#1		read = 32'd2727792933;
		#1		read = 32'd2748439470;
		#1		read = 32'd2769025912;
		#1		read = 32'd2789550200;
		#1		read = 32'd2810010282;
		#1		read = 32'd2830404113;
		#1		read = 32'd2850729651;
		#1		read = 32'd2870984866;
		#1		read = 32'd2891167731;
		#1		read = 32'd2911276228;
		#1		read = 32'd2931308347;
		#1		read = 32'd2951262084;
		#1		read = 32'd2971135444;
		#1		read = 32'd2990926439;
		#1		read = 32'd3010633090;
		#1		read = 32'd3030253428;
		#1		read = 32'd3049785489;
		#1		read = 32'd3069227321;
		#1		read = 32'd3088576979;
		#1		read = 32'd3107832528;
		#1		read = 32'd3126992044;
		#1		read = 32'd3146053609;
		#1		read = 32'd3165015319;
		#1		read = 32'd3183875276;
		#1		read = 32'd3202631595;
		#1		read = 32'd3221282399;
		#1		read = 32'd3239825825;
		#1		read = 32'd3258260018;
		#1		read = 32'd3276583133;
		#1		read = 32'd3294793340;
		#1		read = 32'd3312888817;
		#1		read = 32'd3330867754;
		#1		read = 32'd3348728354;
		#1		read = 32'd3366468830;
		#1		read = 32'd3384087409;
		#1		read = 32'd3401582329;
		#1		read = 32'd3418951839;
		#1		read = 32'd3436194204;
		#1		read = 32'd3453307699;
		#1		read = 32'd3470290613;
		#1		read = 32'd3487141247;
		#1		read = 32'd3503857916;
		#1		read = 32'd3520438949;
		#1		read = 32'd3536882688;
		#1		read = 32'd3553187488;
		#1		read = 32'd3569351718;
		#1		read = 32'd3585373764;
		#1		read = 32'd3601252021;
		#1		read = 32'd3616984902;
		#1		read = 32'd3632570835;
		#1		read = 32'd3648008260;
		#1		read = 32'd3663295635;
		#1		read = 32'd3678431429;
		#1		read = 32'd3693414129;
		#1		read = 32'd3708242238;
		#1		read = 32'd3722914272;
		#1		read = 32'd3737428765;
		#1		read = 32'd3751784264;
		#1		read = 32'd3765979335;
		#1		read = 32'd3780012557;
		#1		read = 32'd3793882528;
		#1		read = 32'd3807587861;
		#1		read = 32'd3821127184;
		#1		read = 32'd3834499145;
		#1		read = 32'd3847702405;
		#1		read = 32'd3860735645;
		#1		read = 32'd3873597561;
		#1		read = 32'd3886286867;
		#1		read = 32'd3898802294;
		#1		read = 32'd3911142591;
		#1		read = 32'd3923306523;
		#1		read = 32'd3935292874;
		#1		read = 32'd3947100447;
		#1		read = 32'd3958728059;
		#1		read = 32'd3970174548;
		#1		read = 32'd3981438769;
		#1		read = 32'd3992519596;
		#1		read = 32'd4003415922;
		#1		read = 32'd4014126655;
		#1		read = 32'd4024650726;
		#1		read = 32'd4034987082;
		#1		read = 32'd4045134689;
		#1		read = 32'd4055092533;
		#1		read = 32'd4064859617;
		#1		read = 32'd4074434965;
		#1		read = 32'd4083817620;
		#1		read = 32'd4093006643;
		#1		read = 32'd4102001115;
		#1		read = 32'd4110800137;
		#1		read = 32'd4119402829;
		#1		read = 32'd4127808331;
		#1		read = 32'd4136015802;
		#1		read = 32'd4144024422;
		#1		read = 32'd4151833389;
		#1		read = 32'd4159441923;
		#1		read = 32'd4166849262;
		#1		read = 32'd4174054667;
		#1		read = 32'd4181057416;
		#1		read = 32'd4187856810;
		#1		read = 32'd4194452168;
		#1		read = 32'd4200842831;
		#1		read = 32'd4207028159;
		#1		read = 32'd4213007535;
		#1		read = 32'd4218780360;
		#1		read = 32'd4224346058;
		#1		read = 32'd4229704070;
		#1		read = 32'd4234853863;
		#1		read = 32'd4239794920;
		#1		read = 32'd4244526748;
		#1		read = 32'd4249048873;
		#1		read = 32'd4253360844;
		#1		read = 32'd4257462228;
		#1		read = 32'd4261352617;
		#1		read = 32'd4265031620;
		#1		read = 32'd4268498870;
		#1		read = 32'd4271754021;
		#1		read = 32'd4274796746;
		#1		read = 32'd4277626742;
		#1		read = 32'd4280243725;
		#1		read = 32'd4282647434;
		#1		read = 32'd4284837628;
		#1		read = 32'd4286814089;
		#1		read = 32'd4288576618;
		#1		read = 32'd4290125040;
		#1		read = 32'd4291459200;
		#1		read = 32'd4292578964;
		#1		read = 32'd4293484220;
		#1		read = 32'd4294174877;
		#1		read = 32'd4294650868;
		#1		read = 32'd4294912143;
		#1		read = 32'd4294958678;
		#1		read = 32'd4294790467;
		#1		read = 32'd4294407527;
		#1		read = 32'd4293809896;
		#1		read = 32'd4292997634;
		#1		read = 32'd4291970823;
		#1		read = 32'd4290729565;
		#1		read = 32'd4289273984;
		#1		read = 32'd4287604226;
		#1		read = 32'd4285720457;
		#1		read = 32'd4283622867;
		#1		read = 32'd4281311665;
		#1		read = 32'd4278787081;
		#1		read = 32'd4276049369;
		#1		read = 32'd4273098802;
		#1		read = 32'd4269935676;
		#1		read = 32'd4266560306;
		#1		read = 32'd4262973030;
		#1		read = 32'd4259174207;
		#1		read = 32'd4255164216;
		#1		read = 32'd4250943459;
		#1		read = 32'd4246512358;
		#1		read = 32'd4241871356;
		#1		read = 32'd4237020917;
		#1		read = 32'd4231961526;
		#1		read = 32'd4226693689;
		#1		read = 32'd4221217933;
		#1		read = 32'd4215534805;
		#1		read = 32'd4209644873;
		#1		read = 32'd4203548727;
		#1		read = 32'd4197246977;
		#1		read = 32'd4190740251;
		#1		read = 32'd4184029202;
		#1		read = 32'd4177114500;
		#1		read = 32'd4169996836;
		#1		read = 32'd4162676923;
		#1		read = 32'd4155155492;
		#1		read = 32'd4147433296;
		#1		read = 32'd4139511106;
		#1		read = 32'd4131389716;
		#1		read = 32'd4123069936;
		#1		read = 32'd4114552599;
		#1		read = 32'd4105838558;
		#1		read = 32'd4096928682;
		#1		read = 32'd4087823863;
		#1		read = 32'd4078525012;
		#1		read = 32'd4069033059;
		#1		read = 32'd4059348952;
		#1		read = 32'd4049473660;
		#1		read = 32'd4039408171;
		#1		read = 32'd4029153490;
		#1		read = 32'd4018710645;
		#1		read = 32'd4008080678;
		#1		read = 32'd3997264653;
		#1		read = 32'd3986263652;
		#1		read = 32'd3975078774;
		#1		read = 32'd3963711138;
		#1		read = 32'd3952161881;
		#1		read = 32'd3940432158;
		#1		read = 32'd3928523141;
		#1		read = 32'd3916436022;
		#1		read = 32'd3904172009;
		#1		read = 32'd3891732328;
		#1		read = 32'd3879118225;
		#1		read = 32'd3866330959;
		#1		read = 32'd3853371810;
		#1		read = 32'd3840242073;
		#1		read = 32'd3826943062;
		#1		read = 32'd3813476107;
		#1		read = 32'd3799842553;
		#1		read = 32'd3786043766;
		#1		read = 32'd3772081123;
		#1		read = 32'd3757956022;
		#1		read = 32'd3743669876;
		#1		read = 32'd3729224111;
		#1		read = 32'd3714620175;
		#1		read = 32'd3699859526;
		#1		read = 32'd3684943640;
		#1		read = 32'd3669874010;
		#1		read = 32'd3654652142;
		#1		read = 32'd3639279559;
		#1		read = 32'd3623757797;
		#1		read = 32'd3608088409;
		#1		read = 32'd3592272961;
		#1		read = 32'd3576313036;
		#1		read = 32'd3560210229;
		#1		read = 32'd3543966151;
		#1		read = 32'd3527582426;
		#1		read = 32'd3511060692;
		#1		read = 32'd3494402601;
		#1		read = 32'd3477609820;
		#1		read = 32'd3460684027;
		#1		read = 32'd3443626915;
		#1		read = 32'd3426440190;
		#1		read = 32'd3409125570;
		#1		read = 32'd3391684787;
		#1		read = 32'd3374119585;
		#1		read = 32'd3356431721;
		#1		read = 32'd3338622963;
		#1		read = 32'd3320695091;
		#1		read = 32'd3302649900;
		#1		read = 32'd3284489193;
		#1		read = 32'd3266214786;
		#1		read = 32'd3247828507;
		#1		read = 32'd3229332195;
		#1		read = 32'd3210727699;
		#1		read = 32'd3192016879;
		#1		read = 32'd3173201606;
		#1		read = 32'd3154283763;
		#1		read = 32'd3135265241;
		#1		read = 32'd3116147941;
		#1		read = 32'd3096933775;
		#1		read = 32'd3077624666;
		#1		read = 32'd3058222543;
		#1		read = 32'd3038729347;
		#1		read = 32'd3019147027;
		#1		read = 32'd2999477541;
		#1		read = 32'd2979722857;
		#1		read = 32'd2959884950;
		#1		read = 32'd2939965803;
		#1		read = 32'd2919967408;
		#1		read = 32'd2899891766;
		#1		read = 32'd2879740884;
		#1		read = 32'd2859516776;
		#1		read = 32'd2839221466;
		#1		read = 32'd2818856983;
		#1		read = 32'd2798425363;
		#1		read = 32'd2777928649;
		#1		read = 32'd2757368891;
		#1		read = 32'd2736748145;
		#1		read = 32'd2716068473;
		#1		read = 32'd2695331944;
		#1		read = 32'd2674540629;
		#1		read = 32'd2653696610;
		#1		read = 32'd2632801970;
		#1		read = 32'd2611858798;
		#1		read = 32'd2590869189;
		#1		read = 32'd2569835242;
		#1		read = 32'd2548759060;
		#1		read = 32'd2527642751;
		#1		read = 32'd2506488427;
		#1		read = 32'd2485298202;
		#1		read = 32'd2464074196;
		#1		read = 32'd2442818531;
		#1		read = 32'd2421533333;
		#1		read = 32'd2400220731;
		#1		read = 32'd2378882854;
		#1		read = 32'd2357521838;
		#1		read = 32'd2336139819;
		#1		read = 32'd2314738934;
		#1		read = 32'd2293321323;
		#1		read = 32'd2271889129;
		#1		read = 32'd2250444495;
		#1		read = 32'd2228989564;
		#1		read = 32'd2207526483;
		#1		read = 32'd2186057398;
		#1		read = 32'd2164584455;
		#1		read = 32'd2143109802;
		#1		read = 32'd2121635587;
		#1		read = 32'd2100163956;
		#1		read = 32'd2078697058;
		#1		read = 32'd2057237038;
		#1		read = 32'd2035786042;
		#1		read = 32'd2014346217;
		#1		read = 32'd1992919704;
		#1		read = 32'd1971508649;
		#1		read = 32'd1950115190;
		#1		read = 32'd1928741468;
		#1		read = 32'd1907389620;
		#1		read = 32'd1886061782;
		#1		read = 32'd1864760085;
		#1		read = 32'd1843486661;
		#1		read = 32'd1822243636;
		#1		read = 32'd1801033134;
		#1		read = 32'd1779857278;
		#1		read = 32'd1758718183;
		#1		read = 32'd1737617965;
		#1		read = 32'd1716558734;
		#1		read = 32'd1695542594;
		#1		read = 32'd1674571648;
		#1		read = 32'd1653647993;
		#1		read = 32'd1632773721;
		#1		read = 32'd1611950920;
		#1		read = 32'd1591181671;
		#1		read = 32'd1570468052;
		#1		read = 32'd1549812134;
		#1		read = 32'd1529215983;
		#1		read = 32'd1508681658;
		#1		read = 32'd1488211213;
		#1		read = 32'd1467806695;
		#1		read = 32'd1447470143;
		#1		read = 32'd1427203593;
		#1		read = 32'd1407009070;
		#1		read = 32'd1386888593;
		#1		read = 32'd1366844176;
		#1		read = 32'd1346877822;
		#1		read = 32'd1326991527;
		#1		read = 32'd1307187281;
		#1		read = 32'd1287467065;
		#1		read = 32'd1267832849;
		#1		read = 32'd1248286597;
		#1		read = 32'd1228830265;
		#1		read = 32'd1209465797;
		#1		read = 32'd1190195130;
		#1		read = 32'd1171020191;
		#1		read = 32'd1151942897;
		#1		read = 32'd1132965157;
		#1		read = 32'd1114088868;
		#1		read = 32'd1095315918;
		#1		read = 32'd1076648183;
		#1		read = 32'd1058087531;
		#1		read = 32'd1039635818;
		#1		read = 32'd1021294888;
		#1		read = 32'd1003066577;
		#1		read = 32'd984952706;
		#1		read = 32'd966955087;
		#1		read = 32'd949075521;
		#1		read = 32'd931315794;
		#1		read = 32'd913677683;
		#1		read = 32'd896162951;
		#1		read = 32'd878773350;
		#1		read = 32'd861510620;
		#1		read = 32'd844376486;
		#1		read = 32'd827372661;
		#1		read = 32'd810500846;
		#1		read = 32'd793762729;
		#1		read = 32'd777159982;
		#1		read = 32'd760694267;
		#1		read = 32'd744367229;
		#1		read = 32'd728180502;
		#1		read = 32'd712135704;
		#1		read = 32'd696234440;
		#1		read = 32'd680478299;
		#1		read = 32'd664868858;
		#1		read = 32'd649407676;
		#1		read = 32'd634096302;
		#1		read = 32'd618936264;
		#1		read = 32'd603929081;
		#1		read = 32'd589076251;
		#1		read = 32'd574379261;
		#1		read = 32'd559839580;
		#1		read = 32'd545458662;
		#1		read = 32'd531237945;
		#1		read = 32'd517178851;
		#1		read = 32'd503282787;
		#1		read = 32'd489551141;
		#1		read = 32'd475985287;
		#1		read = 32'd462586581;
		#1		read = 32'd449356364;
		#1		read = 32'd436295958;
		#1		read = 32'd423406670;
		#1		read = 32'd410689788;
		#1		read = 32'd398146583;
		#1		read = 32'd385778311;
		#1		read = 32'd373586208;
		#1		read = 32'd361571494;
		#1		read = 32'd349735369;
		#1		read = 32'd338079017;
		#1		read = 32'd326603604;
		#1		read = 32'd315310278;
		#1		read = 32'd304200168;
		#1		read = 32'd293274384;
		#1		read = 32'd282534020;
		#1		read = 32'd271980149;
		#1		read = 32'd261613827;
		#1		read = 32'd251436090;
		#1		read = 32'd241447957;
		#1		read = 32'd231650425;
		#1		read = 32'd222044476;
		#1		read = 32'd212631068;
		#1		read = 32'd203411144;
		#1		read = 32'd194385626;
		#1		read = 32'd185555416;
		#1		read = 32'd176921398;
		#1		read = 32'd168484433;
		#1		read = 32'd160245367;
		#1		read = 32'd152205024;
		#1		read = 32'd144364206;
		#1		read = 32'd136723699;
		#1		read = 32'd129284266;
		#1		read = 32'd122046651;
		#1		read = 32'd115011578;
		#1		read = 32'd108179751;
		#1		read = 32'd101551853;
		#1		read = 32'd95128546;
		#1		read = 32'd88910473;
		#1		read = 32'd82898255;
		#1		read = 32'd77092494;
		#1		read = 32'd71493771;
		#1		read = 32'd66102645;
		#1		read = 32'd60919655;
		#1		read = 32'd55945320;
		#1		read = 32'd51180137;
		#1		read = 32'd46624582;
		#1		read = 32'd42279112;
		#1		read = 32'd38144160;
		#1		read = 32'd34220141;
		#1		read = 32'd30507446;
		#1		read = 32'd27006447;
		#1		read = 32'd23717494;
		#1		read = 32'd20640916;
		#1		read = 32'd17777021;
		#1		read = 32'd15126094;
		#1		read = 32'd12688401;
		#1		read = 32'd10464186;
		#1		read = 32'd8453671;
		#1		read = 32'd6657057;
		#1		read = 32'd5074525;
		#1		read = 32'd3706231;
		#1		read = 32'd2552313;
		#1		read = 32'd1612887;
		#1		read = 32'd888046;
		#1		read = 32'd377863;
		#1		read = 32'd82388;
		#1		read = 32'd1652;
		#1		read = 32'd135662;
		#1		read = 32'd484406;
		#1		read = 32'd1047847;
		#1		read = 32'd1825930;
		#1		read = 32'd2818577;
		#1		read = 32'd4025689;
		#1		read = 32'd5447145;
		#1		read = 32'd7082803;
		#1		read = 32'd8932499;
		#1		read = 32'd10996048;
		#1		read = 32'd13273245;
		#1		read = 32'd15763860;
		#1		read = 32'd18467646;
		#1		read = 32'd21384332;
		#1		read = 32'd24513626;
		#1		read = 32'd27855215;
		#1		read = 32'd31408765;
		#1		read = 32'd35173921;
		#1		read = 32'd39150306;
		#1		read = 32'd43337523;
		#1		read = 32'd47735152;
		#1		read = 32'd52342755;
		#1		read = 32'd57159870;
		#1		read = 32'd62186015;
		#1		read = 32'd67420689;
		#1		read = 32'd72863367;
		#1		read = 32'd78513506;
		#1		read = 32'd84370539;
		#1		read = 32'd90433883;
		#1		read = 32'd96702929;
		#1		read = 32'd103177052;
		#1		read = 32'd109855604;
		#1		read = 32'd116737917;
		#1		read = 32'd123823303;
		#1		read = 32'd131111053;
		#1		read = 32'd138600439;
		#1		read = 32'd146290712;
		#1		read = 32'd154181102;
		#1		read = 32'd162270821;
		#1		read = 32'd170559059;
		#1		read = 32'd179044988;
		#1		read = 32'd187727760;
		#1		read = 32'd196606505;
		#1		read = 32'd205680336;
		#1		read = 32'd214948347;
		#1		read = 32'd224409609;
		#1		read = 32'd234063176;
		#1		read = 32'd243908085;
		#1		read = 32'd253943349;
		#1		read = 32'd264167966;
		#1		read = 32'd274580913;
		#1		read = 32'd285181148;
		#1		read = 32'd295967612;
		#1		read = 32'd306939226;
		#1		read = 32'd318094894;
		#1		read = 32'd329433498;
		#1		read = 32'd340953906;
		#1		read = 32'd352654965;
		#1		read = 32'd364535506;
		#1		read = 32'd376594340;
		#1		read = 32'd388830262;
		#1		read = 32'd401242047;
		#1		read = 32'd413828456;
		#1		read = 32'd426588228;
		#1		read = 32'd439520088;
		#1		read = 32'd452622744;
		#1		read = 32'd465894883;
		#1		read = 32'd479335181;
		#1		read = 32'd492942292;
		#1		read = 32'd506714856;
		#1		read = 32'd520651495;
		#1		read = 32'd534750816;
		#1		read = 32'd549011409;
		#1		read = 32'd563431848;
		#1		read = 32'd578010690;
		#1		read = 32'd592746479;
		#1		read = 32'd607637740;
		#1		read = 32'd622682985;
		#1		read = 32'd637880708;
		#1		read = 32'd653229390;
		#1		read = 32'd668727496;
		#1		read = 32'd684373477;
		#1		read = 32'd700165768;
		#1		read = 32'd716102789;
		#1		read = 32'd732182947;
		#1		read = 32'd748404634;
		#1		read = 32'd764766228;
		#1		read = 32'd781266092;
		#1		read = 32'd797902577;
		#1		read = 32'd814674019;
		#1		read = 32'd831578741;
		#1		read = 32'd848615052;
		#1		read = 32'd865781249;
		#1		read = 32'd883075615;
		#1		read = 32'd900496421;
		#1		read = 32'd918041925;
		#1		read = 32'd935710371;
		#1		read = 32'd953499994;
		#1		read = 32'd971409015;
		#1		read = 32'd989435642;
		#1		read = 32'd1007578072;
		#1		read = 32'd1025834493;
		#1		read = 32'd1044203077;
		#1		read = 32'd1062681988;
		#1		read = 32'd1081269379;
		#1		read = 32'd1099963390;
		#1		read = 32'd1118762153;
		#1		read = 32'd1137663786;
		#1		read = 32'd1156666401;
		#1		read = 32'd1175768097;
		#1		read = 32'd1194966963;
		#1		read = 32'd1214261081;
		#1		read = 32'd1233648519;
		#1		read = 32'd1253127341;
		#1		read = 32'd1272695597;
		#1		read = 32'd1292351332;
		#1		read = 32'd1312092579;
		#1		read = 32'd1331917365;
		#1		read = 32'd1351823706;
		#1		read = 32'd1371809613;
		#1		read = 32'd1391873086;
		#1		read = 32'd1412012120;
		#1		read = 32'd1432224701;
		#1		read = 32'd1452508806;
		#1		read = 32'd1472862409;
		#1		read = 32'd1493283473;
		#1		read = 32'd1513769957;
		#1		read = 32'd1534319811;
		#1		read = 32'd1554930982;
		#1		read = 32'd1575601407;
		#1		read = 32'd1596329020;
		#1		read = 32'd1617111748;
		#1		read = 32'd1637947513;
		#1		read = 32'd1658834230;
		#1		read = 32'd1679769813;
		#1		read = 32'd1700752166;
		#1		read = 32'd1721779192;
		#1		read = 32'd1742848789;
		#1		read = 32'd1763958848;
		#1		read = 32'd1785107260;
		#1		read = 32'd1806291909;
		#1		read = 32'd1827510676;
		#1		read = 32'd1848761441;
		#1		read = 32'd1870042078;
		#1		read = 32'd1891350459;
		#1		read = 32'd1912684453;
		#1		read = 32'd1934041926;
		#1		read = 32'd1955420744;
		#1		read = 32'd1976818768;
		#1		read = 32'd1998233858;
		#1		read = 32'd2019663872;
		#1		read = 32'd2041106669;
		#1		read = 32'd2062560104;
		#1		read = 32'd2084022030;
		#1		read = 32'd2105490303;
		#1		read = 32'd2126962775;
		#1		read = 32'd2148437299;
		#1		read = 32'd2169911728;
		#1		read = 32'd2191383914;
		#1		read = 32'd2212851710;
		#1		read = 32'd2234312969;
		#1		read = 32'd2255765546;
		#1		read = 32'd2277207294;
		#1		read = 32'd2298636070;
		#1		read = 32'd2320049731;
		#1		read = 32'd2341446135;
		#1		read = 32'd2362823144;
		#1		read = 32'd2384178618;
		#1		read = 32'd2405510423;
		#1		read = 32'd2426816426;
		#1		read = 32'd2448094496;
		#1		read = 32'd2469342505;
		#1		read = 32'd2490558328;
		#1		read = 32'd2511739844;
		#1		read = 32'd2532884935;
		#1		read = 32'd2553991486;
		#1		read = 32'd2575057387;
		#1		read = 32'd2596080530;
		#1		read = 32'd2617058815;
		#1		read = 32'd2637990142;
		#1		read = 32'd2658872419;
		#1		read = 32'd2679703557;
		#1		read = 32'd2700481474;
		#1		read = 32'd2721204091;
		#1		read = 32'd2741869337;
		#1		read = 32'd2762475145;
		#1		read = 32'd2783019455;
		#1		read = 32'd2803500211;
		#1		read = 32'd2823915366;
		#1		read = 32'd2844262879;
		#1		read = 32'd2864540714;
		#1		read = 32'd2884746844;
		#1		read = 32'd2904879248;
		#1		read = 32'd2924935914;
		#1		read = 32'd2944914834;
		#1		read = 32'd2964814013;
		#1		read = 32'd2984631459;
		#1		read = 32'd3004365191;
		#1		read = 32'd3024013235;
		#1		read = 32'd3043573628;
		#1		read = 32'd3063044412;
		#1		read = 32'd3082423640;
		#1		read = 32'd3101709376;
		#1		read = 32'd3120899690;
		#1		read = 32'd3139992662;
		#1		read = 32'd3158986385;
		#1		read = 32'd3177878959;
		#1		read = 32'd3196668493;
		#1		read = 32'd3215353111;
		#1		read = 32'd3233930942;
		#1		read = 32'd3252400129;
		#1		read = 32'd3270758826;
		#1		read = 32'd3289005195;
		#1		read = 32'd3307137414;
		#1		read = 32'd3325153669;
		#1		read = 32'd3343052157;
		#1		read = 32'd3360831089;
		#1		read = 32'd3378488688;
		#1		read = 32'd3396023187;
		#1		read = 32'd3413432834;
		#1		read = 32'd3430715886;
		#1		read = 32'd3447870616;
		#1		read = 32'd3464895309;
		#1		read = 32'd3481788262;
		#1		read = 32'd3498547785;
		#1		read = 32'd3515172203;
		#1		read = 32'd3531659853;
		#1		read = 32'd3548009087;
		#1		read = 32'd3564218270;
		#1		read = 32'd3580285780;
		#1		read = 32'd3596210011;
		#1		read = 32'd3611989371;
		#1		read = 32'd3627622281;
		#1		read = 32'd3643107179;
		#1		read = 32'd3658442515;
		#1		read = 32'd3673626757;
		#1		read = 32'd3688658386;
		#1		read = 32'd3703535899;
		#1		read = 32'd3718257808;
		#1		read = 32'd3732822641;
		#1		read = 32'd3747228941;
		#1		read = 32'd3761475268;
		#1		read = 32'd3775560197;
		#1		read = 32'd3789482320;
		#1		read = 32'd3803240244;
		#1		read = 32'd3816832594;
		#1		read = 32'd3830258011;
		#1		read = 32'd3843515151;
		#1		read = 32'd3856602690;
		#1		read = 32'd3869519318;
		#1		read = 32'd3882263744;
		#1		read = 32'd3894834694;
		#1		read = 32'd3907230910;
		#1		read = 32'd3919451153;
		#1		read = 32'd3931494200;
		#1		read = 32'd3943358848;
		#1		read = 32'd3955043910;
		#1		read = 32'd3966548217;
		#1		read = 32'd3977870620;
		#1		read = 32'd3989009985;
		#1		read = 32'd3999965199;
		#1		read = 32'd4010735166;
		#1		read = 32'd4021318810;
		#1		read = 32'd4031715072;
		#1		read = 32'd4041922913;
		#1		read = 32'd4051941311;
		#1		read = 32'd4061769264;
		#1		read = 32'd4071405791;
		#1		read = 32'd4080849928;
		#1		read = 32'd4090100729;
		#1		read = 32'd4099157270;
		#1		read = 32'd4108018645;
		#1		read = 32'd4116683969;
		#1		read = 32'd4125152374;
		#1		read = 32'd4133423014;
		#1		read = 32'd4141495062;
		#1		read = 32'd4149367710;
		#1		read = 32'd4157040171;
		#1		read = 32'd4164511679;
		#1		read = 32'd4171781485;
		#1		read = 32'd4178848863;
		#1		read = 32'd4185713107;
		#1		read = 32'd4192373529;
		#1		read = 32'd4198829464;
		#1		read = 32'd4205080266;
		#1		read = 32'd4211125310;
		#1		read = 32'd4216963992;
		#1		read = 32'd4222595727;
		#1		read = 32'd4228019953;
		#1		read = 32'd4233236127;
		#1		read = 32'd4238243727;
		#1		read = 32'd4243042253;
		#1		read = 32'd4247631225;
		#1		read = 32'd4252010184;
		#1		read = 32'd4256178693;
		#1		read = 32'd4260136333;
		#1		read = 32'd4263882710;
		#1		read = 32'd4267417449;
		#1		read = 32'd4270740196;
		#1		read = 32'd4273850619;
		#1		read = 32'd4276748407;
		#1		read = 32'd4279433271;
		#1		read = 32'd4281904941;
		#1		read = 32'd4284163171;
		#1		read = 32'd4286207735;
		#1		read = 32'd4288038429;
		#1		read = 32'd4289655068;
		#1		read = 32'd4291057492;
		#1		read = 32'd4292245561;
		#1		read = 32'd4293219155;
		#1		read = 32'd4293978178;
		#1		read = 32'd4294522552;
		#1		read = 32'd4294852225;
		#1		read = 32'd4294967163;
		#1		read = 32'd4294867354;
		#1		read = 32'd4294552808;
		#1		read = 32'd4294023558;
		#1		read = 32'd4293279655;
		#1		read = 32'd4292321174;
		#1		read = 32'd4291148212;
		#1		read = 32'd4289760884;
		#1		read = 32'd4288159331;
		#1		read = 32'd4286343712;
		#1		read = 32'd4284314209;
		#1		read = 32'd4282071024;
		#1		read = 32'd4279614383;
		#1		read = 32'd4276944530;
		#1		read = 32'd4274061733;
		#1		read = 32'd4270966280;
		#1		read = 32'd4267658480;
		#1		read = 32'd4264138665;
		#1		read = 32'd4260407186;
		#1		read = 32'd4256464416;
		#1		read = 32'd4252310750;
		#1		read = 32'd4247946603;
		#1		read = 32'd4243372412;
		#1		read = 32'd4238588633;
		#1		read = 32'd4233595746;
		#1		read = 32'd4228394249;
		#1		read = 32'd4222984663;
		#1		read = 32'd4217367528;
		#1		read = 32'd4211543407;
		#1		read = 32'd4205512882;
		#1		read = 32'd4199276555;
		#1		read = 32'd4192835051;
		#1		read = 32'd4186189013;
		#1		read = 32'd4179339107;
		#1		read = 32'd4172286016;
		#1		read = 32'd4165030447;
		#1		read = 32'd4157573125;
		#1		read = 32'd4149914796;
		#1		read = 32'd4142056226;
		#1		read = 32'd4133998199;
		#1		read = 32'd4125741523;
		#1		read = 32'd4117287023;
		#1		read = 32'd4108635544;
		#1		read = 32'd4099787952;
		#1		read = 32'd4090745131;
		#1		read = 32'd4081507985;
		#1		read = 32'd4072077438;
		#1		read = 32'd4062454434;
		#1		read = 32'd4052639934;
		#1		read = 32'd4042634920;
		#1		read = 32'd4032440393;
		#1		read = 32'd4022057371;
		#1		read = 32'd4011486894;
		#1		read = 32'd4000730018;
		#1		read = 32'd3989787819;
		#1		read = 32'd3978661391;
		#1		read = 32'd3967351846;
		#1		read = 32'd3955860317;
		#1		read = 32'd3944187951;
		#1		read = 32'd3932335916;
		#1		read = 32'd3920305398;
		#1		read = 32'd3908097598;
		#1		read = 32'd3895713739;
		#1		read = 32'd3883155059;
		#1		read = 32'd3870422812;
		#1		read = 32'd3857518274;
		#1		read = 32'd3844442733;
		#1		read = 32'd3831197497;
		#1		read = 32'd3817783892;
		#1		read = 32'd3804203258;
		#1		read = 32'd3790456953;
		#1		read = 32'd3776546353;
		#1		read = 32'd3762472848;
		#1		read = 32'd3748237845;
		#1		read = 32'd3733842767;
		#1		read = 32'd3719289056;
		#1		read = 32'd3704578165;
		#1		read = 32'd3689711566;
		#1		read = 32'd3674690745;
		#1		read = 32'd3659517205;
		#1		read = 32'd3644192463;
		#1		read = 32'd3628718051;
		#1		read = 32'd3613095518;
		#1		read = 32'd3597326424;
		#1		read = 32'd3581412347;
		#1		read = 32'd3565354878;
		#1		read = 32'd3549155623;
		#1		read = 32'd3532816203;
		#1		read = 32'd3516338250;
		#1		read = 32'd3499723413;
		#1		read = 32'd3482973353;
		#1		read = 32'd3466089745;
		#1		read = 32'd3449074278;
		#1		read = 32'd3431928653;
		#1		read = 32'd3414654584;
		#1		read = 32'd3397253800;
		#1		read = 32'd3379728039;
		#1		read = 32'd3362079055;
		#1		read = 32'd3344308612;
		#1		read = 32'd3326418488;
		#1		read = 32'd3308410471;
		#1		read = 32'd3290286363;
		#1		read = 32'd3272047976;
		#1		read = 32'd3253697132;
		#1		read = 32'd3235235669;
		#1		read = 32'd3216665431;
		#1		read = 32'd3197988276;
		#1		read = 32'd3179206071;
		#1		read = 32'd3160320695;
		#1		read = 32'd3141334036;
		#1		read = 32'd3122247993;
		#1		read = 32'd3103064474;
		#1		read = 32'd3083785398;
		#1		read = 32'd3064412692;
		#1		read = 32'd3044948295;
		#1		read = 32'd3025394151;
		#1		read = 32'd3005752218;
		#1		read = 32'd2986024458;
		#1		read = 32'd2966212845;
		#1		read = 32'd2946319359;
		#1		read = 32'd2926345991;
		#1		read = 32'd2906294737;
		#1		read = 32'd2886167603;
		#1		read = 32'd2865966600;
		#1		read = 32'd2845693750;
		#1		read = 32'd2825351080;
		#1		read = 32'd2804940624;
		#1		read = 32'd2784464422;
		#1		read = 32'd2763924523;
		#1		read = 32'd2743322980;
		#1		read = 32'd2722661854;
		#1		read = 32'd2701943210;
		#1		read = 32'd2681169121;
		#1		read = 32'd2660341664;
		#1		read = 32'd2639462922;
		#1		read = 32'd2618534982;
		#1		read = 32'd2597559937;
		#1		read = 32'd2576539885;
		#1		read = 32'd2555476928;
		#1		read = 32'd2534373171;
		#1		read = 32'd2513230726;
		#1		read = 32'd2492051707;
		#1		read = 32'd2470838231;
		#1		read = 32'd2449592420;
		#1		read = 32'd2428316399;
		#1		read = 32'd2407012294;
		#1		read = 32'd2385682237;
		#1		read = 32'd2364328360;
		#1		read = 32'd2342952798;
		#1		read = 32'd2321557690;
		#1		read = 32'd2300145175;
		#1		read = 32'd2278717394;
		#1		read = 32'd2257276489;
		#1		read = 32'd2235824605;
		#1		read = 32'd2214363888;
		#1		read = 32'd2192896482;
		#1		read = 32'd2171424535;
		#1		read = 32'd2149950194;
		#1		read = 32'd2128475606;
		#1		read = 32'd2107002919;
		#1		read = 32'd2085534280;
		#1		read = 32'd2064071836;
		#1		read = 32'd2042617733;
		#1		read = 32'd2021174117;
		#1		read = 32'd1999743131;
		#1		read = 32'd1978326920;
		#1		read = 32'd1956927624;
		#1		read = 32'd1935547383;
		#1		read = 32'd1914188336;
		#1		read = 32'd1892852618;
		#1		read = 32'd1871542363;
		#1		read = 32'd1850259702;
		#1		read = 32'd1829006763;
		#1		read = 32'd1807785671;
		#1		read = 32'd1786598549;
		#1		read = 32'd1765447516;
		#1		read = 32'd1744334685;
		#1		read = 32'd1723262169;
		#1		read = 32'd1702232075;
		#1		read = 32'd1681246506;
		#1		read = 32'd1660307560;
		#1		read = 32'd1639417331;
		#1		read = 32'd1618577908;
		#1		read = 32'd1597791376;
		#1		read = 32'd1577059812;
		#1		read = 32'd1556385290;
		#1		read = 32'd1535769878;
		#1		read = 32'd1515215636;
		#1		read = 32'd1494724621;
		#1		read = 32'd1474298881;
		#1		read = 32'd1453940459;
		#1		read = 32'd1433651391;
		#1		read = 32'd1413433705;
		#1		read = 32'd1393289424;
		#1		read = 32'd1373220561;
		#1		read = 32'd1353229124;
		#1		read = 32'd1333317112;
		#1		read = 32'd1313486516;
		#1		read = 32'd1293739319;
		#1		read = 32'd1274077496;
		#1		read = 32'd1254503013;
		#1		read = 32'd1235017826;
		#1		read = 32'd1215623886;
		#1		read = 32'd1196323131;
		#1		read = 32'd1177117491;
		#1		read = 32'd1158008887;
		#1		read = 32'd1138999230;
		#1		read = 32'd1120090420;
		#1		read = 32'd1101284349;
		#1		read = 32'd1082582897;
		#1		read = 32'd1063987933;
		#1		read = 32'd1045501319;
		#1		read = 32'd1027124902;
		#1		read = 32'd1008860520;
		#1		read = 32'd990709999;
		#1		read = 32'd972675155;
		#1		read = 32'd954757790;
		#1		read = 32'd936959697;
		#1		read = 32'd919282656;
		#1		read = 32'd901728433;
		#1		read = 32'd884298785;
		#1		read = 32'd866995455;
		#1		read = 32'd849820172;
		#1		read = 32'd832774655;
		#1		read = 32'd815860607;
		#1		read = 32'd799079720;
		#1		read = 32'd782433673;
		#1		read = 32'd765924130;
		#1		read = 32'd749552741;
		#1		read = 32'd733321144;
		#1		read = 32'd717230963;
		#1		read = 32'd701283805;
		#1		read = 32'd685481267;
		#1		read = 32'd669824927;
		#1		read = 32'd654316352;
		#1		read = 32'd638957092;
		#1		read = 32'd623748684;
		#1		read = 32'd608692648;
		#1		read = 32'd593790490;
		#1		read = 32'd579043700;
		#1		read = 32'd564453752;
		#1		read = 32'd550022107;
		#1		read = 32'd535750206;
		#1		read = 32'd521639477;
		#1		read = 32'd507691331;
		#1		read = 32'd493907163;
		#1		read = 32'd480288351;
		#1		read = 32'd466836258;
		#1		read = 32'd453552227;
		#1		read = 32'd440437589;
		#1		read = 32'd427493653;
		#1		read = 32'd414721716;
		#1		read = 32'd402123053;
		#1		read = 32'd389698924;
		#1		read = 32'd377450573;
		#1		read = 32'd365379223;
		#1		read = 32'd353486083;
		#1		read = 32'd341772340;
		#1		read = 32'd330239167;
		#1		read = 32'd318887718;
		#1		read = 32'd307719126;
		#1		read = 32'd296734509;
		#1		read = 32'd285934966;
		#1		read = 32'd275321575;
		#1		read = 32'd264895400;
		#1		read = 32'd254657482;
		#1		read = 32'd244608845;
		#1		read = 32'd234750493;
		#1		read = 32'd225083414;
		#1		read = 32'd215608573;
		#1		read = 32'd206326917;
		#1		read = 32'd197239376;
		#1		read = 32'd188346858;
		#1		read = 32'd179650251;
		#1		read = 32'd171150427;
		#1		read = 32'd162848234;
		#1		read = 32'd154744503;
		#1		read = 32'd146840044;
		#1		read = 32'd139135648;
		#1		read = 32'd131632085;
		#1		read = 32'd124330105;
		#1		read = 32'd117230439;
		#1		read = 32'd110333797;
		#1		read = 32'd103640868;
		#1		read = 32'd97152322;
		#1		read = 32'd90868807;
		#1		read = 32'd84790952;
		#1		read = 32'd78919364;
		#1		read = 32'd73254631;
		#1		read = 32'd67797319;
		#1		read = 32'd62547974;
		#1		read = 32'd57507121;
		#1		read = 32'd52675264;
		#1		read = 32'd48052886;
		#1		read = 32'd43640450;
		#1		read = 32'd39438395;
		#1		read = 32'd35447144;
		#1		read = 32'd31667095;
		#1		read = 32'd28098625;
		#1		read = 32'd24742092;
		#1		read = 32'd21597832;
		#1		read = 32'd18666158;
		#1		read = 32'd15947364;
		#1		read = 32'd13441723;
		#1		read = 32'd11149483;
		#1		read = 32'd9070875;
		#1		read = 32'd7206107;
		#1		read = 32'd5555365;
		#1		read = 32'd4118814;
		#1		read = 32'd2896597;
		#1		read = 32'd1888837;
		#1		read = 32'd1095635;
		#1		read = 32'd517070;
		#1		read = 32'd153200;
		#1		read = 32'd4062;
		#1		read = 32'd69669;
		#1		read = 32'd350016;
		#1		read = 32'd845074;
		#1		read = 32'd1554795;
		#1		read = 32'd2479107;
		#1		read = 32'd3617917;
		#1		read = 32'd4971112;
		#1		read = 32'd6538557;
		#1		read = 32'd8320094;
		#1		read = 32'd10315546;
		#1		read = 32'd12524713;
		#1		read = 32'd14947374;
		#1		read = 32'd17583287;
		#1		read = 32'd20432188;
		#1		read = 32'd23493793;
		#1		read = 32'd26767795;
		#1		read = 32'd30253866;
		#1		read = 32'd33951659;
		#1		read = 32'd37860803;
		#1		read = 32'd41980908;
		#1		read = 32'd46311561;
		#1		read = 32'd50852330;
		#1		read = 32'd55602760;
		#1		read = 32'd60562377;
		#1		read = 32'd65730683;
		#1		read = 32'd71107164;
		#1		read = 32'd76691280;
		#1		read = 32'd82482474;
		#1		read = 32'd88480166;
		#1		read = 32'd94683757;
		#1		read = 32'd101092626;
		#1		read = 32'd107706133;
		#1		read = 32'd114523616;
		#1		read = 32'd121544392;
		#1		read = 32'd128767762;
		#1		read = 32'd136193001;
		#1		read = 32'd143819367;
		#1		read = 32'd151646098;
		#1		read = 32'd159672412;
		#1		read = 32'd167897504;
		#1		read = 32'd176320554;
		#1		read = 32'd184940718;
		#1		read = 32'd193757136;
		#1		read = 32'd202768924;
		#1		read = 32'd211975182;
		#1		read = 32'd221374989;
		#1		read = 32'd230967405;
		#1		read = 32'd240751472;
		#1		read = 32'd250726210;
		#1		read = 32'd260890622;
		#1		read = 32'd271243692;
		#1		read = 32'd281784384;
		#1		read = 32'd292511645;
		#1		read = 32'd303424401;
		#1		read = 32'd314521562;
		#1		read = 32'd325802018;
		#1		read = 32'd337264640;
		#1		read = 32'd348908282;
		#1		read = 32'd360731781;
		#1		read = 32'd372733953;
		#1		read = 32'd384913599;
		#1		read = 32'd397269500;
		#1		read = 32'd409800422;
		#1		read = 32'd422505110;
		#1		read = 32'd435382294;
		#1		read = 32'd448430688;
		#1		read = 32'd461648985;
		#1		read = 32'd475035864;
		#1		read = 32'd488589986;
		#1		read = 32'd502309997;
		#1		read = 32'd516194524;
		#1		read = 32'd530242178;
		#1		read = 32'd544451555;
		#1		read = 32'd558821233;
		#1		read = 32'd573349777;
		#1		read = 32'd588035733;
		#1		read = 32'd602877632;
		#1		read = 32'd617873991;
		#1		read = 32'd633023309;
		#1		read = 32'd648324072;
		#1		read = 32'd663774750;
		#1		read = 32'd679373797;
		#1		read = 32'd695119654;
		#1		read = 32'd711010747;
		#1		read = 32'd727045485;
		#1		read = 32'd743222266;
		#1		read = 32'd759539472;
		#1		read = 32'd775995472;
		#1		read = 32'd792588619;
		#1		read = 32'd809317254;
		#1		read = 32'd826179705;
		#1		read = 32'd843174285;
		#1		read = 32'd860299295;
		#1		read = 32'd877553022;
		#1		read = 32'd894933742;
		#1		read = 32'd912439715;
		#1		read = 32'd930069192;
		#1		read = 32'd947820409;
		#1		read = 32'd965691592;
		#1		read = 32'd983680952;
		#1		read = 32'd1001786692;
		#1		read = 32'd1020007001;
		#1		read = 32'd1038340056;
		#1		read = 32'd1056784025;
		#1		read = 32'd1075337063;
		#1		read = 32'd1093997315;
		#1		read = 32'd1112762914;
		#1		read = 32'd1131631985;
		#1		read = 32'd1150602640;
		#1		read = 32'd1169672982;
		#1		read = 32'd1188841105;
		#1		read = 32'd1208105091;
		#1		read = 32'd1227463014;
		#1		read = 32'd1246912938;
		#1		read = 32'd1266452919;
		#1		read = 32'd1286081002;
		#1		read = 32'd1305795224;
		#1		read = 32'd1325593615;
		#1		read = 32'd1345474194;
		#1		read = 32'd1365434973;
		#1		read = 32'd1385473957;
		#1		read = 32'd1405589141;
		#1		read = 32'd1425778513;
		#1		read = 32'd1446040056;
		#1		read = 32'd1466371742;
		#1		read = 32'd1486771539;
		#1		read = 32'd1507237407;
		#1		read = 32'd1527767298;
		#1		read = 32'd1548359161;
		#1		read = 32'd1569010936;
		#1		read = 32'd1589720558;
		#1		read = 32'd1610485955;
		#1		read = 32'd1631305052;
		#1		read = 32'd1652175766;
		#1		read = 32'd1673096011;
		#1		read = 32'd1694063694;
		#1		read = 32'd1715076718;
		#1		read = 32'd1736132983;
		#1		read = 32'd1757230382;
		#1		read = 32'd1778366807;
		#1		read = 32'd1799540143;
		#1		read = 32'd1820748273;
		#1		read = 32'd1841989076;
		#1		read = 32'd1863260429;
		#1		read = 32'd1884560203;
		#1		read = 32'd1905886270;
		#1		read = 32'd1927236496;
		#1		read = 32'd1948608747;
		#1		read = 32'd1970000885;
		#1		read = 32'd1991410772;
		#1		read = 32'd2012836265;
		#1		read = 32'd2034275223;
		#1		read = 32'd2055725502;
		#1		read = 32'd2077184956;
		#1		read = 32'd2098651440;
		#1		read = 32'd2120122808;
		#1		read = 32'd2141596912;
		#1		read = 32'd2163071604;
		#1		read = 32'd2184544737;
		#1		read = 32'd2206014165;
		#1		read = 32'd2227477739;
		#1		read = 32'd2248933314;
		#1		read = 32'd2270378744;
		#1		read = 32'd2291811885;
		#1		read = 32'd2313230593;
		#1		read = 32'd2334632726;
		#1		read = 32'd2356016145;
		#1		read = 32'd2377378711;
		#1		read = 32'd2398718287;
		#1		read = 32'd2420032740;
		#1		read = 32'd2441319938;
		#1		read = 32'd2462577753;
		#1		read = 32'd2483804059;
		#1		read = 32'd2504996733;
		#1		read = 32'd2526153656;
		#1		read = 32'd2547272713;
		#1		read = 32'd2568351791;
		#1		read = 32'd2589388782;
		#1		read = 32'd2610381583;
		#1		read = 32'd2631328095;
		#1		read = 32'd2652226223;
		#1		read = 32'd2673073877;
		#1		read = 32'd2693868972;
		#1		read = 32'd2714609429;
		#1		read = 32'd2735293174;
		#1		read = 32'd2755918139;
		#1		read = 32'd2776482261;
		#1		read = 32'd2796983483;
		#1		read = 32'd2817419756;
		#1		read = 32'd2837789036;
		#1		read = 32'd2858089286;
		#1		read = 32'd2878318476;
		#1		read = 32'd2898474583;
		#1		read = 32'd2918555592;
		#1		read = 32'd2938559494;
		#1		read = 32'd2958484289;
		#1		read = 32'd2978327985;
		#1		read = 32'd2998088597;
		#1		read = 32'd3017764149;
		#1		read = 32'd3037352674;
		#1		read = 32'd3056852213;
		#1		read = 32'd3076260816;
		#1		read = 32'd3095576541;
		#1		read = 32'd3114797459;
		#1		read = 32'd3133921645;
		#1		read = 32'd3152947189;
		#1		read = 32'd3171872187;
		#1		read = 32'd3190694747;
		#1		read = 32'd3209412987;
		#1		read = 32'd3228025035;
		#1		read = 32'd3246529030;
		#1		read = 32'd3264923121;
		#1		read = 32'd3283205469;
		#1		read = 32'd3301374245;
		#1		read = 32'd3319427634;
		#1		read = 32'd3337363829;
		#1		read = 32'd3355181038;
		#1		read = 32'd3372877477;
		#1		read = 32'd3390451378;
		#1		read = 32'd3407900983;
		#1		read = 32'd3425224548;
		#1		read = 32'd3442420340;
		#1		read = 32'd3459486639;
		#1		read = 32'd3476421739;
		#1		read = 32'd3493223946;
		#1		read = 32'd3509891580;
		#1		read = 32'd3526422975;
		#1		read = 32'd3542816477;
		#1		read = 32'd3559070446;
		#1		read = 32'd3575183259;
		#1		read = 32'd3591153302;
		#1		read = 32'd3606978980;
		#1		read = 32'd3622658709;
		#1		read = 32'd3638190922;
		#1		read = 32'd3653574066;
		#1		read = 32'd3668806601;
		#1		read = 32'd3683887006;
		#1		read = 32'd3698813772;
		#1		read = 32'd3713585406;
		#1		read = 32'd3728200431;
		#1		read = 32'd3742657386;
		#1		read = 32'd3756954825;
		#1		read = 32'd3771091318;
		#1		read = 32'd3785065451;
		#1		read = 32'd3798875828;
		#1		read = 32'd3812521067;
		#1		read = 32'd3825999803;
		#1		read = 32'd3839310689;
		#1		read = 32'd3852452394;
		#1		read = 32'd3865423604;
		#1		read = 32'd3878223021;
		#1		read = 32'd3890849366;
		#1		read = 32'd3903301375;
		#1		read = 32'd3915577804;
		#1		read = 32'd3927677425;
		#1		read = 32'd3939599028;
		#1		read = 32'd3951341421;
		#1		read = 32'd3962903430;
		#1		read = 32'd3974283899;
		#1		read = 32'd3985481689;
		#1		read = 32'd3996495680;
		#1		read = 32'd4007324772;
		#1		read = 32'd4017967882;
		#1		read = 32'd4028423944;
		#1		read = 32'd4038691915;
		#1		read = 32'd4048770765;
		#1		read = 32'd4058659489;
		#1		read = 32'd4068357097;
		#1		read = 32'd4077862619;
		#1		read = 32'd4087175105;
		#1		read = 32'd4096293623;
		#1		read = 32'd4105217262;
		#1		read = 32'd4113945129;
		#1		read = 32'd4122476351;
		#1		read = 32'd4130810076;
		#1		read = 32'd4138945470;
		#1		read = 32'd4146881720;
		#1		read = 32'd4154618031;
		#1		read = 32'd4162153631;
		#1		read = 32'd4169487765;
		#1		read = 32'd4176619700;
		#1		read = 32'd4183548724;
		#1		read = 32'd4190274143;
		#1		read = 32'd4196795284;
		#1		read = 32'd4203111496;
		#1		read = 32'd4209222147;
		#1		read = 32'd4215126626;
		#1		read = 32'd4220824342;
		#1		read = 32'd4226314726;
		#1		read = 32'd4231597228;
		#1		read = 32'd4236671321;
		#1		read = 32'd4241536497;
		#1		read = 32'd4246192269;
		#1		read = 32'd4250638172;
		#1		read = 32'd4254873762;
		#1		read = 32'd4258898614;
		#1		read = 32'd4262712326;
		#1		read = 32'd4266314518;
		#1		read = 32'd4269704828;
		#1		read = 32'd4272882917;
		#1		read = 32'd4275848469;
		#1		read = 32'd4278601186;
		#1		read = 32'd4281140793;
		#1		read = 32'd4283467035;
		#1		read = 32'd4285579682;
		#1		read = 32'd4287478520;
		#1		read = 32'd4289163361;
		#1		read = 32'd4290634036;
		#1		read = 32'd4291890397;
		#1		read = 32'd4292932320;
		#1		read = 32'd4293759699;
		#1		read = 32'd4294372453;
		#1		read = 32'd4294770519;
		#1		read = 32'd4294953859;
		#1		read = 32'd4294922453;
		#1		read = 32'd4294676306;
		#1		read = 32'd4294215440;
		#1		read = 32'd4293539904;
		#1		read = 32'd4292649763;
		#1		read = 32'd4291545108;
		#1		read = 32'd4290226049;
		#1		read = 32'd4288692717;
		#1		read = 32'd4286945265;
		#1		read = 32'd4284983870;
		#1		read = 32'd4282808726;
		#1		read = 32'd4280420052;
		#1		read = 32'd4277818085;
		#1		read = 32'd4275003087;
		#1		read = 32'd4271975339;
		#1		read = 32'd4268735143;
		#1		read = 32'd4265282824;
		#1		read = 32'd4261618727;
		#1		read = 32'd4257743218;
		#1		read = 32'd4253656685;
		#1		read = 32'd4249359536;
		#1		read = 32'd4244852202;
		#1		read = 32'd4240135132;
		#1		read = 32'd4235208799;
		#1		read = 32'd4230073696;
		#1		read = 32'd4224730335;
		#1		read = 32'd4219179251;
		#1		read = 32'd4213420999;
		#1		read = 32'd4207456155;
		#1		read = 32'd4201285316;
		#1		read = 32'd4194909098;
		#1		read = 32'd4188328139;
		#1		read = 32'd4181543098;
		#1		read = 32'd4174554652;
		#1		read = 32'd4167363501;
		#1		read = 32'd4159970364;
		#1		read = 32'd4152375979;
		#1		read = 32'd4144581107;
		#1		read = 32'd4136586527;
		#1		read = 32'd4128393039;
		#1		read = 32'd4120001461;
		#1		read = 32'd4111412633;
		#1		read = 32'd4102627413;
		#1		read = 32'd4093646681;
		#1		read = 32'd4084471335;
		#1		read = 32'd4075102291;
		#1		read = 32'd4065540487;
		#1		read = 32'd4055786878;
		#1		read = 32'd4045842441;
		#1		read = 32'd4035708170;
		#1		read = 32'd4025385078;
		#1		read = 32'd4014874197;
		#1		read = 32'd4004176579;
		#1		read = 32'd3993293293;
		#1		read = 32'd3982225428;
		#1		read = 32'd3970974089;
		#1		read = 32'd3959540404;
		#1		read = 32'd3947925514;
		#1		read = 32'd3936130582;
		#1		read = 32'd3924156786;
		#1		read = 32'd3912005325;
		#1		read = 32'd3899677412;
		#1		read = 32'd3887174282;
		#1		read = 32'd3874497185;
		#1		read = 32'd3861647387;
		#1		read = 32'd3848626174;
		#1		read = 32'd3835434849;
		#1		read = 32'd3822074730;
		#1		read = 32'd3808547153;
		#1		read = 32'd3794853471;
		#1		read = 32'd3780995054;
		#1		read = 32'd3766973287;
		#1		read = 32'd3752789572;
		#1		read = 32'd3738445328;
		#1		read = 32'd3723941989;
		#1		read = 32'd3709281006;
		#1		read = 32'd3694463844;
		#1		read = 32'd3679491985;
		#1		read = 32'd3664366927;
		#1		read = 32'd3649090182;
		#1		read = 32'd3633663277;
		#1		read = 32'd3618087756;
		#1		read = 32'd3602365176;
		#1		read = 32'd3586497108;
		#1		read = 32'd3570485141;
		#1		read = 32'd3554330874;
		#1		read = 32'd3538035924;
		#1		read = 32'd3521601920;
		#1		read = 32'd3505030505;
		#1		read = 32'd3488323336;
		#1		read = 32'd3471482085;
		#1		read = 32'd3454508435;
		#1		read = 32'd3437404084;
		#1		read = 32'd3420170741;
		#1		read = 32'd3402810131;
		#1		read = 32'd3385323990;
		#1		read = 32'd3367714065;
		#1		read = 32'd3349982119;
		#1		read = 32'd3332129923;
		#1		read = 32'd3314159264;
		#1		read = 32'd3296071938;
		#1		read = 32'd3277869755;
		#1		read = 32'd3259554533;
		#1		read = 32'd3241128106;
		#1		read = 32'd3222592315;
		#1		read = 32'd3203949014;
		#1		read = 32'd3185200068;
		#1		read = 32'd3166347350;
		#1		read = 32'd3147392747;
		#1		read = 32'd3128338154;
		#1		read = 32'd3109185477;
		#1		read = 32'd3089936630;
		#1		read = 32'd3070593538;
		#1		read = 32'd3051158137;
		#1		read = 32'd3031632368;
		#1		read = 32'd3012018186;
		#1		read = 32'd2992317551;
		#1		read = 32'd2972532433;
		#1		read = 32'd2952664810;
		#1		read = 32'd2932716671;
		#1		read = 32'd2912690009;
		#1		read = 32'd2892586826;
		#1		read = 32'd2872409135;
		#1		read = 32'd2852158951;
		#1		read = 32'd2831838300;
		#1		read = 32'd2811449214;
		#1		read = 32'd2790993732;
		#1		read = 32'd2770473900;
		#1		read = 32'd2749891770;
		#1		read = 32'd2729249399;
		#1		read = 32'd2708548851;
		#1		read = 32'd2687792198;
		#1		read = 32'd2666981515;
		#1		read = 32'd2646118882;
		#1		read = 32'd2625206386;
		#1		read = 32'd2604246118;
		#1		read = 32'd2583240174;
		#1		read = 32'd2562190655;
		#1		read = 32'd2541099666;
		#1		read = 32'd2519969315;
		#1		read = 32'd2498801716;
		#1		read = 32'd2477598986;
		#1		read = 32'd2456363244;
		#1		read = 32'd2435096615;
		#1		read = 32'd2413801224;
		#1		read = 32'd2392479202;
		#1		read = 32'd2371132681;
		#1		read = 32'd2349763795;
		#1		read = 32'd2328374681;
		#1		read = 32'd2306967478;
		#1		read = 32'd2285544327;
		#1		read = 32'd2264107370;
		#1		read = 32'd2242658750;
		#1		read = 32'd2221200614;
		#1		read = 32'd2199735105;
		#1		read = 32'd2178264372;
		#1		read = 32'd2156790560;
		#1		read = 32'd2135315818;
		#1		read = 32'd2113842293;
		#1		read = 32'd2092372131;
		#1		read = 32'd2070907481;
		#1		read = 32'd2049450488;
		#1		read = 32'd2028003299;
		#1		read = 32'd2006568057;
		#1		read = 32'd1985146907;
		#1		read = 32'd1963741991;
		#1		read = 32'd1942355448;
		#1		read = 32'd1920989418;
		#1		read = 32'd1899646038;
		#1		read = 32'd1878327440;
		#1		read = 32'd1857035759;
		#1		read = 32'd1835773122;
		#1		read = 32'd1814541655;
		#1		read = 32'd1793343483;
		#1		read = 32'd1772180724;
		#1		read = 32'd1751055495;
		#1		read = 32'd1729969909;
		#1		read = 32'd1708926074;
		#1		read = 32'd1687926094;
		#1		read = 32'd1666972070;
		#1		read = 32'd1646066096;
		#1		read = 32'd1625210263;
		#1		read = 32'd1604406658;
		#1		read = 32'd1583657360;
		#1		read = 32'd1562964444;
		#1		read = 32'd1542329979;
		#1		read = 32'd1521756029;
		#1		read = 32'd1501244652;
		#1		read = 32'd1480797898;
		#1		read = 32'd1460417812;
		#1		read = 32'd1440106431;
		#1		read = 32'd1419865788;
		#1		read = 32'd1399697907;
		#1		read = 32'd1379604803;
		#1		read = 32'd1359588486;
		#1		read = 32'd1339650958;
		#1		read = 32'd1319794213;
		#1		read = 32'd1300020236;
		#1		read = 32'd1280331005;
		#1		read = 32'd1260728488;
		#1		read = 32'd1241214646;
		#1		read = 32'd1221791430;
		#1		read = 32'd1202460783;
		#1		read = 32'd1183224637;
		#1		read = 32'd1164084916;
		#1		read = 32'd1145043535;
		#1		read = 32'd1126102396;
		#1		read = 32'd1107263395;
		#1		read = 32'd1088528415;
		#1		read = 32'd1069899329;
		#1		read = 32'd1051378001;
		#1		read = 32'd1032966283;
		#1		read = 32'd1014666016;
		#1		read = 32'd996479029;
		#1		read = 32'd978407142;
		#1		read = 32'd960452161;
		#1		read = 32'd942615883;
		#1		read = 32'd924900090;
		#1		read = 32'd907306555;
		#1		read = 32'd889837037;
		#1		read = 32'd872493282;
		#1		read = 32'd855277025;
		#1		read = 32'd838189988;
		#1		read = 32'd821233878;
		#1		read = 32'd804410393;
		#1		read = 32'd787721214;
		#1		read = 32'd771168010;
		#1		read = 32'd754752437;
		#1		read = 32'd738476135;
		#1		read = 32'd722340733;
		#1		read = 32'd706347845;
		#1		read = 32'd690499068;
		#1		read = 32'd674795989;
		#1		read = 32'd659240177;
		#1		read = 32'd643833189;
		#1		read = 32'd628576564;
		#1		read = 32'd613471829;
		#1		read = 32'd598520493;
		#1		read = 32'd583724053;
		#1		read = 32'd569083987;
		#1		read = 32'd554601760;
		#1		read = 32'd540278820;
		#1		read = 32'd526116599;
		#1		read = 32'd512116513;
		#1		read = 32'd498279962;
		#1		read = 32'd484608331;
		#1		read = 32'd471102986;
		#1		read = 32'd457765277;
		#1		read = 32'd444596539;
		#1		read = 32'd431598088;
		#1		read = 32'd418771224;
		#1		read = 32'd406117231;
		#1		read = 32'd393637372;
		#1		read = 32'd381332896;
		#1		read = 32'd369205034;
		#1		read = 32'd357254999;
		#1		read = 32'd345483984;
		#1		read = 32'd333893169;
		#1		read = 32'd322483710;
		#1		read = 32'd311256751;
		#1		read = 32'd300213412;
		#1		read = 32'd289354799;
		#1		read = 32'd278681997;
		#1		read = 32'd268196074;
		#1		read = 32'd257898078;
		#1		read = 32'd247789039;
		#1		read = 32'd237869968;
		#1		read = 32'd228141857;
		#1		read = 32'd218605678;
		#1		read = 32'd209262385;
		#1		read = 32'd200112913;
		#1		read = 32'd191158177;
		#1		read = 32'd182399071;
		#1		read = 32'd173836472;
		#1		read = 32'd165471236;
		#1		read = 32'd157304200;
		#1		read = 32'd149336180;
		#1		read = 32'd141567974;
		#1		read = 32'd134000357;
		#1		read = 32'd126634086;
		#1		read = 32'd119469899;
		#1		read = 32'd112508512;
		#1		read = 32'd105750620;
		#1		read = 32'd99196901;
		#1		read = 32'd92848008;
		#1		read = 32'd86704577;
		#1		read = 32'd80767222;
		#1		read = 32'd75036537;
		#1		read = 32'd69513095;
		#1		read = 32'd64197448;
		#1		read = 32'd59090128;
		#1		read = 32'd54191646;
		#1		read = 32'd49502491;
		#1		read = 32'd45023133;
		#1		read = 32'd40754019;
		#1		read = 32'd36695576;
		#1		read = 32'd32848210;
		#1		read = 32'd29212306;
		#1		read = 32'd25788228;
		#1		read = 32'd22576317;
		#1		read = 32'd19576895;
		#1		read = 32'd16790262;
		#1		read = 32'd14216696;
		#1		read = 32'd11856456;
		#1		read = 32'd9709776;
		#1		read = 32'd7776872;
		#1		read = 32'd6057937;
		#1		read = 32'd4553143;
		#1		read = 32'd3262640;
		#1		read = 32'd2186557;
		#1		read = 32'd1325002;
		#1		read = 32'd678062;
		#1		read = 32'd245800;
		#1		read = 32'd28260;
		#1		read = 32'd25464;
		#1		read = 32'd237411;
		#1		read = 32'd664082;
		#1		read = 32'd1305433;
		#1		read = 32'd2161400;
		#1		read = 32'd3231897;
		#1		read = 32'd4516818;
		#1		read = 32'd6016033;
		#1		read = 32'd7729394;
		#1		read = 32'd9656728;
		#1		read = 32'd11797843;
		#1		read = 32'd14152525;
		#1		read = 32'd16720538;
		#1		read = 32'd19501626;
		#1		read = 32'd22495510;
		#1		read = 32'd25701892;
		#1		read = 32'd29120449;
		#1		read = 32'd32750841;
		#1		read = 32'd36592705;
		#1		read = 32'd40645656;
		#1		read = 32'd44909289;
		#1		read = 32'd49383178;
		#1		read = 32'd54066875;
		#1		read = 32'd58959912;
		#1		read = 32'd64061800;
		#1		read = 32'd69372028;
		#1		read = 32'd74890066;
		#1		read = 32'd80615361;
		#1		read = 32'd86547341;
		#1		read = 32'd92685413;
		#1		read = 32'd99028963;
		#1		read = 32'd105577358;
		#1		read = 32'd112329941;
		#1		read = 32'd119286037;
		#1		read = 32'd126444952;
		#1		read = 32'd133805969;
		#1		read = 32'd141368352;
		#1		read = 32'd149131345;
		#1		read = 32'd157094171;
		#1		read = 32'd165256035;
		#1		read = 32'd173616120;
		#1		read = 32'd182173590;
		#1		read = 32'd190927589;
		#1		read = 32'd199877242;
		#1		read = 32'd209021655;
		#1		read = 32'd218359911;
		#1		read = 32'd227891079;
		#1		read = 32'd237614204;
		#1		read = 32'd247528315;
		#1		read = 32'd257632420;
		#1		read = 32'd267925508;
		#1		read = 32'd278406550;
		#1		read = 32'd289074499;
		#1		read = 32'd299928287;
		#1		read = 32'd310966829;
		#1		read = 32'd322189021;
		#1		read = 32'd333593741;
		#1		read = 32'd345179848;
		#1		read = 32'd356946185;
		#1		read = 32'd368891573;
		#1		read = 32'd381014820;
		#1		read = 32'd393314711;
		#1		read = 32'd405790018;
		#1		read = 32'd418439494;
		#1		read = 32'd431261872;
		#1		read = 32'd444255870;
		#1		read = 32'd457420191;
		#1		read = 32'd470753516;
		#1		read = 32'd484254513;
		#1		read = 32'd497921831;
		#1		read = 32'd511754104;
		#1		read = 32'd525749949;
		#1		read = 32'd539907965;
		#1		read = 32'd554226738;
		#1		read = 32'd568704835;
		#1		read = 32'd583340809;
		#1		read = 32'd598133196;
		#1		read = 32'd613080517;
		#1		read = 32'd628181276;
		#1		read = 32'd643433965;
		#1		read = 32'd658837057;
		#1		read = 32'd674389013;
		#1		read = 32'd690088277;
		#1		read = 32'd705933279;
		#1		read = 32'd721922435;
		#1		read = 32'd738054146;
		#1		read = 32'd754326799;
		#1		read = 32'd770738766;
		#1		read = 32'd787288407;
		#1		read = 32'd803974066;
		#1		read = 32'd820794075;
		#1		read = 32'd837746752;
		#1		read = 32'd854830401;
		#1		read = 32'd872043315;
		#1		read = 32'd889383771;
		#1		read = 32'd906850037;
		#1		read = 32'd924440365;
		#1		read = 32'd942152996;
		#1		read = 32'd959986159;
		#1		read = 32'd977938071;
		#1		read = 32'd996006937;
		#1		read = 32'd1014190949;
		#1		read = 32'd1032488289;
		#1		read = 32'd1050897129;
		#1		read = 32'd1069415626;
		#1		read = 32'd1088041928;
		#1		read = 32'd1106774175;
		#1		read = 32'd1125610491;
		#1		read = 32'd1144548993;
		#1		read = 32'd1163587789;
		#1		read = 32'd1182724973;
		#1		read = 32'd1201958632;
		#1		read = 32'd1221286843;
		#1		read = 32'd1240707673;
		#1		read = 32'd1260219179;
		#1		read = 32'd1279819411;
		#1		read = 32'd1299506410;
		#1		read = 32'd1319278205;
		#1		read = 32'd1339132819;
		#1		read = 32'd1359068269;
		#1		read = 32'd1379082559;
		#1		read = 32'd1399173689;
		#1		read = 32'd1419339649;
		#1		read = 32'd1439578422;
		#1		read = 32'd1459887986;
		#1		read = 32'd1480266309;
		#1		read = 32'd1500711353;
		#1		read = 32'd1521221073;
		#1		read = 32'd1541793420;
		#1		read = 32'd1562426334;
		#1		read = 32'd1583117755;
		#1		read = 32'd1603865611;
		#1		read = 32'd1624667828;
		#1		read = 32'd1645522327;
		#1		read = 32'd1666427021;
		#1		read = 32'd1687379821;
		#1		read = 32'd1708378631;
		#1		read = 32'd1729421351;
		#1		read = 32'd1750505876;
		#1		read = 32'd1771630100;
		#1		read = 32'd1792791908;
		#1		read = 32'd1813989185;
		#1		read = 32'd1835219811;
		#1		read = 32'd1856481663;
		#1		read = 32'd1877772616;
		#1		read = 32'd1899090539;
		#1		read = 32'd1920433301;
		#1		read = 32'd1941798768;
		#1		read = 32'd1963184804;
		#1		read = 32'd1984589269;
		#1		read = 32'd2006010024;
		#1		read = 32'd2027444925;
		#1		read = 32'd2048891831;
		#1		read = 32'd2070348595;
		#1		read = 32'd2091813073;
		#1		read = 32'd2113283118;
		#1		read = 32'd2134756584;
		#1		read = 32'd2156231321;
		#1		read = 32'd2177705184;
		#1		read = 32'd2199176025;
		#1		read = 32'd2220641697;
		#1		read = 32'd2242100053;
		#1		read = 32'd2263548947;
		#1		read = 32'd2284986235;
		#1		read = 32'd2306409773;
		#1		read = 32'd2327817418;
		#1		read = 32'd2349207031;
		#1		read = 32'd2370576470;
		#1		read = 32'd2391923601;
		#1		read = 32'd2413246288;
		#1		read = 32'd2434542399;
		#1		read = 32'd2455809805;
		#1		read = 32'd2477046378;
		#1		read = 32'd2498249995;
		#1		read = 32'd2519418535;
		#1		read = 32'd2540549883;
		#1		read = 32'd2561641924;
		#1		read = 32'd2582692550;
		#1		read = 32'd2603699655;
		#1		read = 32'd2624661139;
		#1		read = 32'd2645574906;
		#1		read = 32'd2666438864;
		#1		read = 32'd2687250926;
		#1		read = 32'd2708009013;
		#1		read = 32'd2728711047;
		#1		read = 32'd2749354960;
		#1		read = 32'd2769938685;
		#1		read = 32'd2790460166;
		#1		read = 32'd2810917349;
		#1		read = 32'd2831308190;
		#1		read = 32'd2851630649;
		#1		read = 32'd2871882693;
		#1		read = 32'd2892062299;
		#1		read = 32'd2912167447;
		#1		read = 32'd2932196127;
		#1		read = 32'd2952146337;
		#1		read = 32'd2972016081;
		#1		read = 32'd2991803373;
		#1		read = 32'd3011506233;
		#1		read = 32'd3031122692;
		#1		read = 32'd3050650788;
		#1		read = 32'd3070088567;
		#1		read = 32'd3089434087;
		#1		read = 32'd3108685413;
		#1		read = 32'd3127840619;
		#1		read = 32'd3146897791;
		#1		read = 32'd3165855022;
		#1		read = 32'd3184710416;
		#1		read = 32'd3203462089;
		#1		read = 32'd3222108165;
		#1		read = 32'd3240646779;
		#1		read = 32'd3259076078;
		#1		read = 32'd3277394219;
		#1		read = 32'd3295599369;
		#1		read = 32'd3313689709;
		#1		read = 32'd3331663429;
		#1		read = 32'd3349518732;
		#1		read = 32'd3367253833;
		#1		read = 32'd3384866958;
		#1		read = 32'd3402356345;
		#1		read = 32'd3419720246;
		#1		read = 32'd3436956925;
		#1		read = 32'd3454064657;
		#1		read = 32'd3471041732;
		#1		read = 32'd3487886453;
		#1		read = 32'd3504597134;
		#1		read = 32'd3521172105;
		#1		read = 32'd3537609709;
		#1		read = 32'd3553908301;
		#1		read = 32'd3570066252;
		#1		read = 32'd3586081945;
		#1		read = 32'd3601953780;
		#1		read = 32'd3617680170;
		#1		read = 32'd3633259540;
		#1		read = 32'd3648690335;
		#1		read = 32'd3663971010;
		#1		read = 32'd3679100038;
		#1		read = 32'd3694075905;
		#1		read = 32'd3708897114;
		#1		read = 32'd3723562183;
		#1		read = 32'd3738069646;
		#1		read = 32'd3752418051;
		#1		read = 32'd3766605965;
		#1		read = 32'd3780631967;
		#1		read = 32'd3794494656;
		#1		read = 32'd3808192645;
		#1		read = 32'd3821724565;
		#1		read = 32'd3835089062;
		#1		read = 32'd3848284800;
		#1		read = 32'd3861310459;
		#1		read = 32'd3874164737;
		#1		read = 32'd3886846348;
		#1		read = 32'd3899354025;
		#1		read = 32'd3911686516;
		#1		read = 32'd3923842588;
		#1		read = 32'd3935821025;
		#1		read = 32'd3947620631;
		#1		read = 32'd3959240224;
		#1		read = 32'd3970678643;
		#1		read = 32'd3981934744;
		#1		read = 32'd3993007402;
		#1		read = 32'd4003895508;
		#1		read = 32'd4014597975;
		#1		read = 32'd4025113732;
		#1		read = 32'd4035441728;
		#1		read = 32'd4045580930;
		#1		read = 32'd4055530323;
		#1		read = 32'd4065288913;
		#1		read = 32'd4074855724;
		#1		read = 32'd4084229800;
		#1		read = 32'd4093410203;
		#1		read = 32'd4102396014;
		#1		read = 32'd4111186336;
		#1		read = 32'd4119780290;
		#1		read = 32'd4128177015;
		#1		read = 32'd4136375673;
		#1		read = 32'd4144375443;
		#1		read = 32'd4152175526;
		#1		read = 32'd4159775141;
		#1		read = 32'd4167173529;
		#1		read = 32'd4174369949;
		#1		read = 32'd4181363682;
		#1		read = 32'd4188154030;
		#1		read = 32'd4194740311;
		#1		read = 32'd4201121869;
		#1		read = 32'd4207298065;
		#1		read = 32'd4213268281;
		#1		read = 32'd4219031920;
		#1		read = 32'd4224588406;
		#1		read = 32'd4229937184;
		#1		read = 32'd4235077717;
		#1		read = 32'd4240009493;
		#1		read = 32'd4244732019;
		#1		read = 32'd4249244821;
		#1		read = 32'd4253547449;
		#1		read = 32'd4257639472;
		#1		read = 32'd4261520481;
		#1		read = 32'd4265190089;
		#1		read = 32'd4268647927;
		#1		read = 32'd4271893651;
		#1		read = 32'd4274926936;
		#1		read = 32'd4277747478;
		#1		read = 32'd4280354995;
		#1		read = 32'd4282749228;
		#1		read = 32'd4284929935;
		#1		read = 32'd4286896899;
		#1		read = 32'd4288649924;
		#1		read = 32'd4290188835;
		#1		read = 32'd4291513476;
		#1		read = 32'd4292623716;
		#1		read = 32'd4293519444;
		#1		read = 32'd4294200570;
		#1		read = 32'd4294667027;
		#1		read = 32'd4294918766;
		#1		read = 32'd4294955764;
		#1		read = 32'd4294778017;
		#1		read = 32'd4294385542;
		#1		read = 32'd4293778379;
		#1		read = 32'd4292956587;
		#1		read = 32'd4291920251;
		#1		read = 32'd4290669472;
		#1		read = 32'd4289204377;
		#1		read = 32'd4287525111;
		#1		read = 32'd4285631843;
		#1		read = 32'd4283524762;
		#1		read = 32'd4281204079;
		#1		read = 32'd4278670025;
		#1		read = 32'd4275922855;
		#1		read = 32'd4272962842;
		#1		read = 32'd4269790284;
		#1		read = 32'd4266405496;
		#1		read = 32'd4262808818;
		#1		read = 32'd4259000609;
		#1		read = 32'd4254981250;
		#1		read = 32'd4250751144;
		#1		read = 32'd4246310712;
		#1		read = 32'd4241660399;
		#1		read = 32'd4236800671;
		#1		read = 32'd4231732012;
		#1		read = 32'd4226454930;
		#1		read = 32'd4220969953;
		#1		read = 32'd4215277629;
		#1		read = 32'd4209378527;
		#1		read = 32'd4203273238;
		#1		read = 32'd4196962371;
		#1		read = 32'd4190446558;
		#1		read = 32'd4183726451;
		#1		read = 32'd4176802721;
		#1		read = 32'd4169676061;
		#1		read = 32'd4162347183;
		#1		read = 32'd4154816820;
		#1		read = 32'd4147085726;
		#1		read = 32'd4139154674;
		#1		read = 32'd4131024456;
		#1		read = 32'd4122695885;
		#1		read = 32'd4114169795;
		#1		read = 32'd4105447038;
		#1		read = 32'd4096528486;
		#1		read = 32'd4087415031;
		#1		read = 32'd4078107585;
		#1		read = 32'd4068607078;
		#1		read = 32'd4058914461;
		#1		read = 32'd4049030701;
		#1		read = 32'd4038956789;
		#1		read = 32'd4028693731;
		#1		read = 32'd4018242553;
		#1		read = 32'd4007604302;
		#1		read = 32'd3996780039;
		#1		read = 32'd3985770849;
		#1		read = 32'd3974577831;
		#1		read = 32'd3963202106;
		#1		read = 32'd3951644810;
		#1		read = 32'd3939907099;
		#1		read = 32'd3927990148;
		#1		read = 32'd3915895148;
		#1		read = 32'd3903623307;
		#1		read = 32'd3891175855;
		#1		read = 32'd3878554034;
		#1		read = 32'd3865759108;
		#1		read = 32'd3852792356;
		#1		read = 32'd3839655075;
		#1		read = 32'd3826348577;
		#1		read = 32'd3812874195;
		#1		read = 32'd3799233275;
		#1		read = 32'd3785427181;
		#1		read = 32'd3771457295;
		#1		read = 32'd3757325012;
		#1		read = 32'd3743031746;
		#1		read = 32'd3728578927;
		#1		read = 32'd3713968000;
		#1		read = 32'd3699200426;
		#1		read = 32'd3684277681;
		#1		read = 32'd3669201259;
		#1		read = 32'd3653972665;
		#1		read = 32'd3638593424;
		#1		read = 32'd3623065074;
		#1		read = 32'd3607389166;
		#1		read = 32'd3591567269;
		#1		read = 32'd3575600965;
		#1		read = 32'd3559491850;
		#1		read = 32'd3543241536;
		#1		read = 32'd3526851647;
		#1		read = 32'd3510323823;
		#1		read = 32'd3493659715;
		#1		read = 32'd3476860992;
		#1		read = 32'd3459929331;
		#1		read = 32'd3442866427;
		#1		read = 32'd3425673986;
		#1		read = 32'd3408353727;
		#1		read = 32'd3390907382;
		#1		read = 32'd3373336695;
		#1		read = 32'd3355643424;
		#1		read = 32'd3337829339;
		#1		read = 32'd3319896219;
		#1		read = 32'd3301845860;
		#1		read = 32'd3283680065;
		#1		read = 32'd3265400651;
		#1		read = 32'd3247009447;
		#1		read = 32'd3228508291;
		#1		read = 32'd3209899034;
		#1		read = 32'd3191183535;
		#1		read = 32'd3172363668;
		#1		read = 32'd3153441314;
		#1		read = 32'd3134418364;
		#1		read = 32'd3115296722;
		#1		read = 32'd3096078300;
		#1		read = 32'd3076765019;
		#1		read = 32'd3057358810;
		#1		read = 32'd3037861615;
		#1		read = 32'd3018275382;
		#1		read = 32'd2998602071;
		#1		read = 32'd2978843650;
		#1		read = 32'd2959002092;
		#1		read = 32'd2939079384;
		#1		read = 32'd2919077517;
		#1		read = 32'd2898998490;
		#1		read = 32'd2878844313;
		#1		read = 32'd2858617001;
		#1		read = 32'd2838318576;
		#1		read = 32'd2817951068;
		#1		read = 32'd2797516514;
		#1		read = 32'd2777016957;
		#1		read = 32'd2756454447;
		#1		read = 32'd2735831040;
		#1		read = 32'd2715148800;
		#1		read = 32'd2694409793;
		#1		read = 32'd2673616094;
		#1		read = 32'd2652769783;
		#1		read = 32'd2631872943;
		#1		read = 32'd2610927665;
		#1		read = 32'd2589936042;
		#1		read = 32'd2568900175;
		#1		read = 32'd2547822167;
		#1		read = 32'd2526704124;
		#1		read = 32'd2505548161;
		#1		read = 32'd2484356391;
		#1		read = 32'd2463130934;
		#1		read = 32'd2441873912;
		#1		read = 32'd2420587452;
		#1		read = 32'd2399273682;
		#1		read = 32'd2377934733;
		#1		read = 32'd2356572739;
		#1		read = 32'd2335189836;
		#1		read = 32'd2313788163;
		#1		read = 32'd2292369859;
		#1		read = 32'd2270937067;
		#1		read = 32'd2249491930;
		#1		read = 32'd2228036592;
		#1		read = 32'd2206573199;
		#1		read = 32'd2185103896;
		#1		read = 32'd2163630832;
		#1		read = 32'd2142156153;
		#1		read = 32'd2120682007;
		#1		read = 32'd2099210541;
		#1		read = 32'd2077743903;
		#1		read = 32'd2056284238;
		#1		read = 32'd2034833693;
		#1		read = 32'd2013394413;
		#1		read = 32'd1991968542;
		#1		read = 32'd1970558222;
		#1		read = 32'd1949165594;
		#1		read = 32'd1927792799;
		#1		read = 32'd1906441972;
		#1		read = 32'd1885115249;
		#1		read = 32'd1863814763;
		#1		read = 32'd1842542643;
		#1		read = 32'd1821301017;
		#1		read = 32'd1800092009;
		#1		read = 32'd1778917740;
		#1		read = 32'd1757780328;
		#1		read = 32'd1736681885;
		#1		read = 32'd1715624522;
		#1		read = 32'd1694610345;
		#1		read = 32'd1673641455;
		#1		read = 32'd1652719948;
		#1		read = 32'd1631847918;
		#1		read = 32'd1611027450;
		#1		read = 32'd1590260628;
		#1		read = 32'd1569549528;
		#1		read = 32'd1548896220;
		#1		read = 32'd1528302771;
		#1		read = 32'd1507771239;
		#1		read = 32'd1487303679;
		#1		read = 32'd1466902135;
		#1		read = 32'd1446568649;
		#1		read = 32'd1426305254;
		#1		read = 32'd1406113977;
		#1		read = 32'd1385996835;
		#1		read = 32'd1365955842;
		#1		read = 32'd1345993001;
		#1		read = 32'd1326110308;
		#1		read = 32'd1306309752;
		#1		read = 32'd1286593312;
		#1		read = 32'd1266962961;
		#1		read = 32'd1247420661;
		#1		read = 32'd1227968367;
		#1		read = 32'd1208608023;
		#1		read = 32'd1189341567;
		#1		read = 32'd1170170923;
		#1		read = 32'd1151098010;
		#1		read = 32'd1132124735;
		#1		read = 32'd1113252995;
		#1		read = 32'd1094484677;
		#1		read = 32'd1075821659;
		#1		read = 32'd1057265805;
		#1		read = 32'd1038818972;
		#1		read = 32'd1020483005;
		#1		read = 32'd1002259737;
		#1		read = 32'd984150991;
		#1		read = 32'd966158576;
		#1		read = 32'd948284294;
		#1		read = 32'd930529930;
		#1		read = 32'd912897260;
		#1		read = 32'd895388048;
		#1		read = 32'd878004045;
		#1		read = 32'd860746989;
		#1		read = 32'd843618605;
		#1		read = 32'd826620606;
		#1		read = 32'd809754693;
		#1		read = 32'd793022552;
		#1		read = 32'd776425855;
		#1		read = 32'd759966263;
		#1		read = 32'd743645422;
		#1		read = 32'd727464964;
		#1		read = 32'd711426506;
		#1		read = 32'd695531652;
		#1		read = 32'd679781993;
		#1		read = 32'd664179103;
		#1		read = 32'd648724541;
		#1		read = 32'd633419855;
		#1		read = 32'd618266573;
		#1		read = 32'd603266212;
		#1		read = 32'd588420272;
		#1		read = 32'd573730236;
		#1		read = 32'd559197575;
		#1		read = 32'd544823740;
		#1		read = 32'd530610171;
		#1		read = 32'd516558287;
		#1		read = 32'd502669495;
		#1		read = 32'd488945183;
		#1		read = 32'd475386723;
		#1		read = 32'd461995471;
		#1		read = 32'd448772767;
		#1		read = 32'd435719933;
		#1		read = 32'd422838273;
		#1		read = 32'd410129077;
		#1		read = 32'd397593614;
		#1		read = 32'd385233139;
		#1		read = 32'd373048888;
		#1		read = 32'd361042079;
		#1		read = 32'd349213912;
		#1		read = 32'd337565571;
		#1		read = 32'd326098220;
		#1		read = 32'd314813006;
		#1		read = 32'd303711058;
		#1		read = 32'd292793485;
		#1		read = 32'd282061380;
		#1		read = 32'd271515816;
		#1		read = 32'd261157847;
		#1		read = 32'd250988508;
		#1		read = 32'd241008818;
		#1		read = 32'd231219774;
		#1		read = 32'd221622354;
		#1		read = 32'd212217519;
		#1		read = 32'd203006209;
		#1		read = 32'd193989345;
		#1		read = 32'd185167829;
		#1		read = 32'd176542543;
		#1		read = 32'd168114349;
		#1		read = 32'd159884091;
		#1		read = 32'd151852590;
		#1		read = 32'd144020652;
		#1		read = 32'd136389058;
		#1		read = 32'd128958571;
		#1		read = 32'd121729936;
		#1		read = 32'd114703874;
		#1		read = 32'd107881089;
		#1		read = 32'd101262262;
		#1		read = 32'd94848055;
		#1		read = 32'd88639111;
		#1		read = 32'd82636049;
		#1		read = 32'd76839470;
		#1		read = 32'd71249954;
		#1		read = 32'd65868059;
		#1		read = 32'd60694324;
		#1		read = 32'd55729267;
		#1		read = 32'd50973383;
		#1		read = 32'd46427148;
		#1		read = 32'd42091018;
		#1		read = 32'd37965425;
		#1		read = 32'd34050782;
		#1		read = 32'd30347480;
		#1		read = 32'd26855890;
		#1		read = 32'd23576362;
		#1		read = 32'd20509222;
		#1		read = 32'd17654778;
		#1		read = 32'd15013315;
		#1		read = 32'd12585097;
		#1		read = 32'd10370368;
		#1		read = 32'd8369347;
		#1		read = 32'd6582237;
		#1		read = 32'd5009215;
		#1		read = 32'd3650439;
		#1		read = 32'd2506044;
		#1		read = 32'd1576145;
		#1		read = 32'd860835;
		#1		read = 32'd360185;
		#1		read = 32'd74246;
		#1		read = 32'd3047;
		#1		read = 32'd146593;
		#1		read = 32'd504872;
		#1		read = 32'd1077846;
		#1		read = 32'd1865460;
		#1		read = 32'd2867633;
		#1		read = 32'd4084266;
		#1		read = 32'd5515237;
		#1		read = 32'd7160404;
		#1		read = 32'd9019601;
		#1		read = 32'd11092642;
		#1		read = 32'd13379321;
		#1		read = 32'd15879409;
		#1		read = 32'd18592655;
		#1		read = 32'd21518788;
		#1		read = 32'd24657516;
		#1		read = 32'd28008526;
		#1		read = 32'd31571480;
		#1		read = 32'd35346025;
		#1		read = 32'd39331781;
		#1		read = 32'd43528350;
		#1		read = 32'd47935314;
		#1		read = 32'd52552230;
		#1		read = 32'd57378638;
		#1		read = 32'd62414055;
		#1		read = 32'd67657977;
		#1		read = 32'd73109880;
		#1		read = 32'd78769218;
		#1		read = 32'd84635426;
		#1		read = 32'd90707917;
		#1		read = 32'd96986085;
		#1		read = 32'd103469300;
		#1		read = 32'd110156915;
		#1		read = 32'd117048260;
		#1		read = 32'd124142648;
		#1		read = 32'd131439368;
		#1		read = 32'd138937691;
		#1		read = 32'd146636867;
		#1		read = 32'd154536126;
		#1		read = 32'd162634677;
		#1		read = 32'd170931713;
		#1		read = 32'd179426401;
		#1		read = 32'd188117894;
		#1		read = 32'd197005322;
		#1		read = 32'd206087795;
		#1		read = 32'd215364407;
		#1		read = 32'd224834230;
		#1		read = 32'd234496315;
		#1		read = 32'd244349698;
		#1		read = 32'd254393392;
		#1		read = 32'd264626394;
		#1		read = 32'd275047680;
		#1		read = 32'd285656208;
		#1		read = 32'd296450917;
		#1		read = 32'd307430729;
		#1		read = 32'd318594543;
		#1		read = 32'd329941245;
		#1		read = 32'd341469700;
		#1		read = 32'd353178755;
		#1		read = 32'd365067239;
		#1		read = 32'd377133963;
		#1		read = 32'd389377720;
		#1		read = 32'd401797287;
		#1		read = 32'd414391421;
		#1		read = 32'd427158862;
		#1		read = 32'd440098335;
		#1		read = 32'd453208544;
		#1		read = 32'd466488180;
		#1		read = 32'd479935914;
		#1		read = 32'd493550401;
		#1		read = 32'd507330281;
		#1		read = 32'd521274174;
		#1		read = 32'd535380687;
		#1		read = 32'd549648408;
		#1		read = 32'd564075912;
		#1		read = 32'd578661756;
		#1		read = 32'd593404480;
		#1		read = 32'd608302611;
		#1		read = 32'd623354659;
		#1		read = 32'd638559118;
		#1		read = 32'd653914468;
		#1		read = 32'd669419175;
		#1		read = 32'd685071686;
		#1		read = 32'd700870438;
		#1		read = 32'd716813849;
		#1		read = 32'd732900326;
		#1		read = 32'd749128261;
		#1		read = 32'd765496030;
		#1		read = 32'd782001996;
		#1		read = 32'd798644510;
		#1		read = 32'd815421906;
		#1		read = 32'd832332507;
		#1		read = 32'd849374623;
		#1		read = 32'd866546548;
		#1		read = 32'd883846566;
		#1		read = 32'd901272946;
		#1		read = 32'd918823947;
		#1		read = 32'd936497812;
		#1		read = 32'd954292775;
		#1		read = 32'd972207056;
		#1		read = 32'd990238864;
		#1		read = 32'd1008386395;
		#1		read = 32'd1026647835;
		#1		read = 32'd1045021358;
		#1		read = 32'd1063505126;
		#1		read = 32'd1082097291;
		#1		read = 32'd1100795994;
		#1		read = 32'd1119599365;
		#1		read = 32'd1138505523;
		#1		read = 32'd1157512578;
		#1		read = 32'd1176618630;
		#1		read = 32'd1195821767;
		#1		read = 32'd1215120069;
		#1		read = 32'd1234511607;
		#1		read = 32'd1253994442;
		#1		read = 32'd1273566625;
		#1		read = 32'd1293226198;
		#1		read = 32'd1312971197;
		#1		read = 32'd1332799646;
		#1		read = 32'd1352709564;
		#1		read = 32'd1372698957;
		#1		read = 32'd1392765829;
		#1		read = 32'd1412908172;
		#1		read = 32'd1433123971;
		#1		read = 32'd1453411206;
		#1		read = 32'd1473767848;
		#1		read = 32'd1494191861;
		#1		read = 32'd1514681202;
		#1		read = 32'd1535233823;
		#1		read = 32'd1555847669;
		#1		read = 32'd1576520678;
		#1		read = 32'd1597250782;
		#1		read = 32'd1618035909;
		#1		read = 32'd1638873981;
		#1		read = 32'd1659762913;
		#1		read = 32'd1680700617;
		#1		read = 32'd1701684999;
		#1		read = 32'd1722713960;
		#1		read = 32'd1743785398;
		#1		read = 32'd1764897205;
		#1		read = 32'd1786047271;
		#1		read = 32'd1807233480;
		#1		read = 32'd1828453714;
		#1		read = 32'd1849705850;
		#1		read = 32'd1870987764;
		#1		read = 32'd1892297328;
		#1		read = 32'd1913632410;
		#1		read = 32'd1934990876;
		#1		read = 32'd1956370592;
		#1		read = 32'd1977769419;
		#1		read = 32'd1999185218;
		#1		read = 32'd2020615846;
		#1		read = 32'd2042059160;
		#1		read = 32'd2063513017;
		#1		read = 32'd2084975271;
		#1		read = 32'd2106443776;
		#1		read = 32'd2127916385;
		#1		read = 32'd2149390950;
		#1		read = 32'd2170865325;
		#1		read = 32'd2192337362;
		#1		read = 32'd2213804913;
		#1		read = 32'd2235265832;
		#1		read = 32'd2256717973;
		#1		read = 32'd2278159191;
		#1		read = 32'd2299587341;
		#1		read = 32'd2321000281;
		#1		read = 32'd2342395869;
		#1		read = 32'd2363771967;
		#1		read = 32'd2385126436;
		#1		read = 32'd2406457140;
		#1		read = 32'd2427761948;
		#1		read = 32'd2449038728;
		#1		read = 32'd2470285353;
		#1		read = 32'd2491499697;
		#1		read = 32'd2512679641;
		#1		read = 32'd2533823065;
		#1		read = 32'd2554927856;
		#1		read = 32'd2575991902;
		#1		read = 32'd2597013098;
		#1		read = 32'd2617989342;
		#1		read = 32'd2638918535;
		#1		read = 32'd2659798585;
		#1		read = 32'd2680627404;
		#1		read = 32'd2701402909;
		#1		read = 32'd2722123023;
		#1		read = 32'd2742785673;
		#1		read = 32'd2763388794;
		#1		read = 32'd2783930325;
		#1		read = 32'd2804408211;
		#1		read = 32'd2824820406;
		#1		read = 32'd2845164867;
		#1		read = 32'd2865439561;
		#1		read = 32'd2885642460;
		#1		read = 32'd2905771543;
		#1		read = 32'd2925824799;
		#1		read = 32'd2945800221;
		#1		read = 32'd2965695812;
		#1		read = 32'd2985509582;
		#1		read = 32'd3005239551;
		#1		read = 32'd3024883744;
		#1		read = 32'd3044440199;
		#1		read = 32'd3063906958;
		#1		read = 32'd3083282076;
		#1		read = 32'd3102563615;
		#1		read = 32'd3121749647;
		#1		read = 32'd3140838253;
		#1		read = 32'd3159827524;
		#1		read = 32'd3178715562;
		#1		read = 32'd3197500477;
		#1		read = 32'd3216180392;
		#1		read = 32'd3234753437;
		#1		read = 32'd3253217757;
		#1		read = 32'd3271571504;
		#1		read = 32'd3289812844;
		#1		read = 32'd3307939951;
		#1		read = 32'd3325951014;
		#1		read = 32'd3343844231;
		#1		read = 32'd3361617813;
		#1		read = 32'd3379269982;
		#1		read = 32'd3396798974;
		#1		read = 32'd3414203036;
		#1		read = 32'd3431480426;
		#1		read = 32'd3448629418;
		#1		read = 32'd3465648297;
		#1		read = 32'd3482535360;
		#1		read = 32'd3499288919;
		#1		read = 32'd3515907298;
		#1		read = 32'd3532388837;
		#1		read = 32'd3548731886;
		#1		read = 32'd3564934811;
		#1		read = 32'd3580995992;
		#1		read = 32'd3596913824;
		#1		read = 32'd3612686713;
		#1		read = 32'd3628313084;
		#1		read = 32'd3643791373;
		#1		read = 32'd3659120032;
		#1		read = 32'd3674297529;
		#1		read = 32'd3689322346;
		#1		read = 32'd3704192980;
		#1		read = 32'd3718907944;
		#1		read = 32'd3733465768;
		#1		read = 32'd3747864994;
		#1		read = 32'd3762104184;
		#1		read = 32'd3776181913;
		#1		read = 32'd3790096774;
		#1		read = 32'd3803847374;
		#1		read = 32'd3817432340;
		#1		read = 32'd3830850312;
		#1		read = 32'd3844099949;
		#1		read = 32'd3857179926;
		#1		read = 32'd3870088934;
		#1		read = 32'd3882825683;
		#1		read = 32'd3895388900;
		#1		read = 32'd3907777328;
		#1		read = 32'd3919989727;
		#1		read = 32'd3932024878;
		#1		read = 32'd3943881576;
		#1		read = 32'd3955558635;
		#1		read = 32'd3967054889;
		#1		read = 32'd3978369187;
		#1		read = 32'd3989500398;
		#1		read = 32'd4000447409;
		#1		read = 32'd4011209125;
		#1		read = 32'd4021784470;
		#1		read = 32'd4032172386;
		#1		read = 32'd4042371835;
		#1		read = 32'd4052381797;
		#1		read = 32'd4062201271;
		#1		read = 32'd4071829274;
		#1		read = 32'd4081264845;
		#1		read = 32'd4090507039;
		#1		read = 32'd4099554932;
		#1		read = 32'd4108407620;
		#1		read = 32'd4117064217;
		#1		read = 32'd4125523858;
		#1		read = 32'd4133785696;
		#1		read = 32'd4141848906;
		#1		read = 32'd4149712681;
		#1		read = 32'd4157376234;
		#1		read = 32'd4164838800;
		#1		read = 32'd4172099633;
		#1		read = 32'd4179158005;
		#1		read = 32'd4186013212;
		#1		read = 32'd4192664567;
		#1		read = 32'd4199111406;
		#1		read = 32'd4205353084;
		#1		read = 32'd4211388976;
		#1		read = 32'd4217218480;
		#1		read = 32'd4222841012;
		#1		read = 32'd4228256010;
		#1		read = 32'd4233462933;
		#1		read = 32'd4238461259;
		#1		read = 32'd4243250489;
		#1		read = 32'd4247830145;
		#1		read = 32'd4252199767;
		#1		read = 32'd4256358920;
		#1		read = 32'd4260307187;
		#1		read = 32'd4264044173;
		#1		read = 32'd4267569505;
		#1		read = 32'd4270882830;
		#1		read = 32'd4273983817;
		#1		read = 32'd4276872156;
		#1		read = 32'd4279547558;
		#1		read = 32'd4282009755;
		#1		read = 32'd4284258501;
		#1		read = 32'd4286293572;
		#1		read = 32'd4288114763;
		#1		read = 32'd4289721893;
		#1		read = 32'd4291114801;
		#1		read = 32'd4292293348;
		#1		read = 32'd4293257415;
		#1		read = 32'd4294006907;
		#1		read = 32'd4294541748;
		#1		read = 32'd4294861886;
		#1		read = 32'd4294967287;
		#1		read = 32'd4294857942;
		#1		read = 32'd4294533861;
		#1		read = 32'd4293995077;
		#1		read = 32'd4293241643;
		#1		read = 32'd4292273636;
		#1		read = 32'd4291091151;
		#1		read = 32'd4289694307;
		#1		read = 32'd4288083244;
		#1		read = 32'd4286258123;
		#1		read = 32'd4284219126;
		#1		read = 32'd4281966458;
		#1		read = 32'd4279500342;
		#1		read = 32'd4276821027;
		#1		read = 32'd4273928780;
		#1		read = 32'd4270823891;
		#1		read = 32'd4267506669;
		#1		read = 32'd4263977446;
		#1		read = 32'd4260236576;
		#1		read = 32'd4256284433;
		#1		read = 32'd4252121411;
		#1		read = 32'd4247747927;
		#1		read = 32'd4243164418;
		#1		read = 32'd4238371343;
		#1		read = 32'd4233369181;
		#1		read = 32'd4228158432;
		#1		read = 32'd4222739618;
		#1		read = 32'd4217113279;
		#1		read = 32'd4211279980;
		#1		read = 32'd4205240302;
		#1		read = 32'd4198994850;
		#1		read = 32'd4192544249;
		#1		read = 32'd4185889144;
		#1		read = 32'd4179030200;
		#1		read = 32'd4171968103;
		#1		read = 32'd4164703559;
		#1		read = 32'd4157237295;
		#1		read = 32'd4149570057;
		#1		read = 32'd4141702612;
		#1		read = 32'd4133635747;
		#1		read = 32'd4125370268;
		#1		read = 32'd4116907003;
		#1		read = 32'd4108246796;
		#1		read = 32'd4099390515;
		#1		read = 32'd4090339045;
		#1		read = 32'd4081093291;
		#1		read = 32'd4071654178;
		#1		read = 32'd4062022649;
		#1		read = 32'd4052199668;
		#1		read = 32'd4042186217;
		#1		read = 32'd4031983297;
		#1		read = 32'd4021591929;
		#1		read = 32'd4011013151;
		#1		read = 32'd4000248022;
		#1		read = 32'd3989297619;
		#1		read = 32'd3978163035;
		#1		read = 32'd3966845385;
		#1		read = 32'd3955345800;
		#1		read = 32'd3943665431;
		#1		read = 32'd3931805445;
		#1		read = 32'd3919767028;
		#1		read = 32'd3907551384;
		#1		read = 32'd3895159735;
		#1		read = 32'd3882593320;
		#1		read = 32'd3869853396;
		#1		read = 32'd3856941236;
		#1		read = 32'd3843858131;
		#1		read = 32'd3830605391;
		#1		read = 32'd3817184339;
		#1		read = 32'd3803596319;
		#1		read = 32'd3789842689;
		#1		read = 32'd3775924825;
		#1		read = 32'd3761844118;
		#1		read = 32'd3747601976;
		#1		read = 32'd3733199824;
		#1		read = 32'd3718639101;
		#1		read = 32'd3703921264;
		#1		read = 32'd3689047785;
		#1		read = 32'd3674020150;
		#1		read = 32'd3658839863;
		#1		read = 32'd3643508442;
		#1		read = 32'd3628027420;
		#1		read = 32'd3612398344;
		#1		read = 32'd3596622778;
		#1		read = 32'd3580702300;
		#1		read = 32'd3564638500;
		#1		read = 32'd3548432987;
		#1		read = 32'd3532087380;
		#1		read = 32'd3515603313;
		#1		read = 32'd3498982436;
		#1		read = 32'd3482226410;
		#1		read = 32'd3465336910;
		#1		read = 32'd3448315627;
		#1		read = 32'd3431164261;
		#1		read = 32'd3413884529;
		#1		read = 32'd3396478157;
		#1		read = 32'd3378946887;
		#1		read = 32'd3361292472;
		#1		read = 32'd3343516677;
		#1		read = 32'd3325621279;
		#1		read = 32'd3307608069;
		#1		read = 32'd3289478847;
		#1		read = 32'd3271235427;
		#1		read = 32'd3252879632;
		#1		read = 32'd3234413299;
		#1		read = 32'd3215838273;
		#1		read = 32'd3197156414;
		#1		read = 32'd3178369587;
		#1		read = 32'd3159479673;
		#1		read = 32'd3140488561;
		#1		read = 32'd3121398148;
		#1		read = 32'd3102210345;
		#1		read = 32'd3082927070;
		#1		read = 32'd3063550251;
		#1		read = 32'd3044081827;
		#1		read = 32'd3024523744;
		#1		read = 32'd3004877957;
		#1		read = 32'd2985146431;
		#1		read = 32'd2965331140;
		#1		read = 32'd2945434065;
		#1		read = 32'd2925457196;
		#1		read = 32'd2905402529;
		#1		read = 32'd2885272072;
		#1		read = 32'd2865067836;
		#1		read = 32'd2844791843;
		#1		read = 32'd2824446119;
		#1		read = 32'd2804032700;
		#1		read = 32'd2783553626;
		#1		read = 32'd2763010945;
		#1		read = 32'd2742406713;
		#1		read = 32'd2721742989;
		#1		read = 32'd2701021839;
		#1		read = 32'd2680245336;
		#1		read = 32'd2659415557;
		#1		read = 32'd2638534585;
		#1		read = 32'd2617604509;
		#1		read = 32'd2596627421;
		#1		read = 32'd2575605419;
		#1		read = 32'd2554540605;
		#1		read = 32'd2533435086;
		#1		read = 32'd2512290972;
		#1		read = 32'd2491110378;
		#1		read = 32'd2469895421;
		#1		read = 32'd2448648223;
		#1		read = 32'd2427370909;
		#1		read = 32'd2406065607;
		#1		read = 32'd2384734447;
		#1		read = 32'd2363379561;
		#1		read = 32'd2342003087;
		#1		read = 32'd2320607160;
		#1		read = 32'd2299193922;
		#1		read = 32'd2277765512;
		#1		read = 32'd2256324074;
		#1		read = 32'd2234871753;
		#1		read = 32'd2213410692;
		#1		read = 32'd2191943039;
		#1		read = 32'd2170470941;
		#1		read = 32'd2148996543;
		#1		read = 32'd2127521994;
		#1		read = 32'd2106049441;
		#1		read = 32'd2084581032;
		#1		read = 32'd2063118913;
		#1		read = 32'd2041665230;
		#1		read = 32'd2020222129;
		#1		read = 32'd1998791754;
		#1		read = 32'd1977376248;
		#1		read = 32'd1955977753;
		#1		read = 32'd1934598408;
		#1		read = 32'd1913240352;
		#1		read = 32'd1891905719;
		#1		read = 32'd1870596645;
		#1		read = 32'd1849315258;
		#1		read = 32'd1828063689;
		#1		read = 32'd1806844061;
		#1		read = 32'd1785658496;
		#1		read = 32'd1764509114;
		#1		read = 32'd1743398029;
		#1		read = 32'd1722327352;
		#1		read = 32'd1701299191;
		#1		read = 32'd1680315648;
		#1		read = 32'd1659378821;
		#1		read = 32'd1638490804;
		#1		read = 32'd1617653686;
		#1		read = 32'd1596869550;
		#1		read = 32'd1576140476;
		#1		read = 32'd1555468535;
		#1		read = 32'd1534855795;
		#1		read = 32'd1514304318;
		#1		read = 32'd1493816158;
		#1		read = 32'd1473393364;
		#1		read = 32'd1453037979;
		#1		read = 32'd1432752037;
		#1		read = 32'd1412537569;
		#1		read = 32'd1392396594;
		#1		read = 32'd1372331127;
		#1		read = 32'd1352343175;
		#1		read = 32'd1332434736;
		#1		read = 32'd1312607802;
		#1		read = 32'd1292864354;
		#1		read = 32'd1273206368;
		#1		read = 32'd1253635808;
		#1		read = 32'd1234154633;
		#1		read = 32'd1214764790;
		#1		read = 32'd1195468218;
		#1		read = 32'd1176266846;
		#1		read = 32'd1157162596;
		#1		read = 32'd1138157377;
		#1		read = 32'd1119253089;
		#1		read = 32'd1100451624;
		#1		read = 32'd1081754861;
		#1		read = 32'd1063164670;
		#1		read = 32'd1044682910;
		#1		read = 32'd1026311429;
		#1		read = 32'd1008052065;
		#1		read = 32'd989906643;
		#1		read = 32'd971876977;
		#1		read = 32'd953964871;
		#1		read = 32'd936172116;
		#1		read = 32'd918500492;
		#1		read = 32'd900951764;
		#1		read = 32'd883527689;
		#1		read = 32'd866230008;
		#1		read = 32'd849060451;
		#1		read = 32'd832020736;
		#1		read = 32'd815112566;
		#1		read = 32'd798337632;
		#1		read = 32'd781697611;
		#1		read = 32'd765194168;
		#1		read = 32'd748828953;
		#1		read = 32'd732603602;
		#1		read = 32'd716519737;
		#1		read = 32'd700578968;
		#1		read = 32'd684782889;
		#1		read = 32'd669133078;
		#1		read = 32'd653631101;
		#1		read = 32'd638278508;
		#1		read = 32'd623076834;
		#1		read = 32'd608027599;
		#1		read = 32'd593132309;
		#1		read = 32'd578392453;
		#1		read = 32'd563809505;
		#1		read = 32'd549384922;
		#1		read = 32'd535120148;
		#1		read = 32'd521016610;
		#1		read = 32'd507075716;
		#1		read = 32'd493298862;
		#1		read = 32'd479687425;
		#1		read = 32'd466242767;
		#1		read = 32'd452966231;
		#1		read = 32'd439859145;
		#1		read = 32'd426922820;
		#1		read = 32'd414158550;
		#1		read = 32'd401567611;
		#1		read = 32'd389151263;
		#1		read = 32'd376910746;
		#1		read = 32'd364847284;
		#1		read = 32'd352962085;
		#1		read = 32'd341256337;
		#1		read = 32'd329731210;
		#1		read = 32'd318387856;
		#1		read = 32'd307227411;
		#1		read = 32'd296250990;
		#1		read = 32'd285459690;
		#1		read = 32'd274854591;
		#1		read = 32'd264436754;
		#1		read = 32'd254207220;
		#1		read = 32'd244167012;
		#1		read = 32'd234317134;
		#1		read = 32'd224658570;
		#1		read = 32'd215192288;
		#1		read = 32'd205919234;
		#1		read = 32'd196840334;
		#1		read = 32'd187956497;
		#1		read = 32'd179268611;
		#1		read = 32'd170777545;
		#1		read = 32'd162484147;
		#1		read = 32'd154389249;
		#1		read = 32'd146493658;
		#1		read = 32'd138798164;
		#1		read = 32'd131303537;
		#1		read = 32'd124010526;
		#1		read = 32'd116919861;
		#1		read = 32'd110032251;
		#1		read = 32'd103348384;
		#1		read = 32'd96868929;
		#1		read = 32'd90594534;
		#1		read = 32'd84525826;
		#1		read = 32'd78663412;
		#1		read = 32'd73007878;
		#1		read = 32'd67559791;
		#1		read = 32'd62319693;
		#1		read = 32'd57288111;
		#1		read = 32'd52465546;
		#1		read = 32'd47852482;
		#1		read = 32'd43449378;
		#1		read = 32'd39256677;
		#1		read = 32'd35274796;
		#1		read = 32'd31504135;
		#1		read = 32'd27945069;
		#1		read = 32'd24597956;
		#1		read = 32'd21463129;
		#1		read = 32'd18540903;
		#1		read = 32'd15831570;
		#1		read = 32'd13335399;
		#1		read = 32'd11052642;
		#1		read = 32'd8983526;
		#1		read = 32'd7128259;
		#1		read = 32'd5487025;
		#1		read = 32'd4059989;
		#1		read = 32'd2847293;
		#1		read = 32'd1849060;
		#1		read = 32'd1065388;
		#1		read = 32'd496356;
		#1		read = 32'd142021;
		#1		read = 32'd2419;
		#1		read = 32'd77562;
		#1		read = 32'd367445;
		#1		read = 32'd872037;
		#1		read = 32'd1591289;
		#1		read = 32'd2525128;
		#1		read = 32'd3673462;
		#1		read = 32'd5036174;
		#1		read = 32'd6613130;
		#1		read = 32'd8404171;
		#1		read = 32'd10409117;
		#1		read = 32'd12627770;
		#1		read = 32'd15059907;
		#1		read = 32'd17705284;
		#1		read = 32'd20563637;
		#1		read = 32'd23634680;
		#1		read = 32'd26918106;
		#1		read = 32'd30413588;
		#1		read = 32'd34120774;
		#1		read = 32'd38039295;
		#1		read = 32'd42168759;
		#1		read = 32'd46508752;
		#1		read = 32'd51058841;
		#1		read = 32'd55818571;
		#1		read = 32'd60787466;
		#1		read = 32'd65965028;
		#1		read = 32'd71350741;
		#1		read = 32'd76944065;
		#1		read = 32'd82744442;
		#1		read = 32'd88751290;
		#1		read = 32'd94964010;
		#1		read = 32'd101381981;
		#1		read = 32'd108004560;
		#1		read = 32'd114831085;
		#1		read = 32'd121860873;
		#1		read = 32'd129093223;
		#1		read = 32'd136527409;
		#1		read = 32'd144162690;
		#1		read = 32'd151998301;
		#1		read = 32'd160033459;
		#1		read = 32'd168267360;
		#1		read = 32'd176699181;
		#1		read = 32'd185328079;
		#1		read = 32'd194153191;
		#1		read = 32'd203173634;
		#1		read = 32'd212388507;
		#1		read = 32'd221796888;
		#1		read = 32'd231397835;
		#1		read = 32'd241190390;
		#1		read = 32'd251173572;
		#1		read = 32'd261346384;
		#1		read = 32'd271707808;
		#1		read = 32'd282256808;
		#1		read = 32'd292992329;
		#1		read = 32'd303913298;
		#1		read = 32'd315018622;
		#1		read = 32'd326307191;
		#1		read = 32'd337777877;
		#1		read = 32'd349429531;
		#1		read = 32'd361260989;
		#1		read = 32'd373271068;
		#1		read = 32'd385458567;
		#1		read = 32'd397822267;
		#1		read = 32'd410360932;
		#1		read = 32'd423073307;
		#1		read = 32'd435958122;
		#1		read = 32'd449014088;
		#1		read = 32'd462239900;
		#1		read = 32'd475634235;
		#1		read = 32'd489195753;
		#1		read = 32'd502923098;
		#1		read = 32'd516814899;
		#1		read = 32'd530869765;
		#1		read = 32'd545086290;
		#1		read = 32'd559463055;
		#1		read = 32'd573998620;
		#1		read = 32'd588691532;
		#1		read = 32'd603540322;
		#1		read = 32'd618543505;
		#1		read = 32'd633699581;
		#1		read = 32'd649007034;
		#1		read = 32'd664464333;
		#1		read = 32'd680069933;
		#1		read = 32'd695822274;
		#1		read = 32'd711719779;
		#1		read = 32'd727760859;
		#1		read = 32'd743943911;
		#1		read = 32'd760267315;
		#1		read = 32'd776729440;
		#1		read = 32'd793328639;
		#1		read = 32'd810063252;
		#1		read = 32'd826931607;
		#1		read = 32'd843932015;
		#1		read = 32'd861062778;
		#1		read = 32'd878322181;
		#1		read = 32'd895708500;
		#1		read = 32'd913219995;
		#1		read = 32'd930854915;
		#1		read = 32'd948611498;
		#1		read = 32'd966487966;
		#1		read = 32'd984482533;
		#1		read = 32'd1002593399;
		#1		read = 32'd1020818754;
		#1		read = 32'd1039156774;
		#1		read = 32'd1057605625;
		#1		read = 32'd1076163464;
		#1		read = 32'd1094828433;
		#1		read = 32'd1113598668;
		#1		read = 32'd1132472290;
		#1		read = 32'd1151447412;
		#1		read = 32'd1170522137;
		#1		read = 32'd1189694557;
		#1		read = 32'd1208962756;
		#1		read = 32'd1228324805;
		#1		read = 32'd1247778770;
		#1		read = 32'd1267322705;
		#1		read = 32'd1286954655;
		#1		read = 32'd1306672657;
		#1		read = 32'd1326474739;
		#1		read = 32'd1346358922;
		#1		read = 32'd1366323217;
		#1		read = 32'd1386365627;
		#1		read = 32'd1406484148;
		#1		read = 32'd1426676768;
		#1		read = 32'd1446941469;
		#1		read = 32'd1467276223;
		#1		read = 32'd1487678997;
		#1		read = 32'd1508147752;
		#1		read = 32'd1528680439;
		#1		read = 32'd1549275006;
		#1		read = 32'd1569929394;
		#1		read = 32'd1590641536;
		#1		read = 32'd1611409362;
		#1		read = 32'd1632230796;
		#1		read = 32'd1653103754;
		#1		read = 32'd1674026149;
		#1		read = 32'd1694995890;
		#1		read = 32'd1716010879;
		#1		read = 32'd1737069016;
		#1		read = 32'd1758168193;
		#1		read = 32'd1779306302;
		#1		read = 32'd1800481228;
		#1		read = 32'd1821690854;
		#1		read = 32'd1842933059;
		#1		read = 32'd1864205719;
		#1		read = 32'd1885506706;
		#1		read = 32'd1906833891;
		#1		read = 32'd1928185141;
		#1		read = 32'd1949558320;
		#1		read = 32'd1970951291;
		#1		read = 32'd1992361916;
		#1		read = 32'd2013788053;
		#1		read = 32'd2035227559;
		#1		read = 32'd2056678291;
		#1		read = 32'd2078138103;
		#1		read = 32'd2099604850;
		#1		read = 32'd2121076384;
		#1		read = 32'd2142550560;
		#1		read = 32'd2164025228;
		#1		read = 32'd2185498243;
		#1		read = 32'd2206967456;
		#1		read = 32'd2228430720;
		#1		read = 32'd2249885890;
		#1		read = 32'd2271330820;
		#1		read = 32'd2292763366;
		#1		read = 32'd2314181383;
		#1		read = 32'd2335582731;
		#1		read = 32'd2356965269;
		#1		read = 32'd2378326859;
		#1		read = 32'd2399665365;
		#1		read = 32'd2420978653;
		#1		read = 32'd2442264591;
		#1		read = 32'd2463521052;
		#1		read = 32'd2484745909;
		#1		read = 32'd2505937041;
		#1		read = 32'd2527092327;
		#1		read = 32'd2548209653;
		#1		read = 32'd2569286907;
		#1		read = 32'd2590321980;
		#1		read = 32'd2611312770;
		#1		read = 32'd2632257178;
		#1		read = 32'd2653153109;
		#1		read = 32'd2673998473;
		#1		read = 32'd2694791186;
		#1		read = 32'd2715529168;
		#1		read = 32'd2736210347;
		#1		read = 32'd2756832654;
		#1		read = 32'd2777394026;
		#1		read = 32'd2797892407;
		#1		read = 32'd2818325749;
		#1		read = 32'd2838692006;
		#1		read = 32'd2858989144;
		#1		read = 32'd2879215131;
		#1		read = 32'd2899367946;
		#1		read = 32'd2919445573;
		#1		read = 32'd2939446005;
		#1		read = 32'd2959367240;
		#1		read = 32'd2979207289;
		#1		read = 32'd2998964165;
		#1		read = 32'd3018635895;
		#1		read = 32'd3038220509;
		#1		read = 32'd3057716051;
		#1		read = 32'd3077120570;
		#1		read = 32'd3096432127;
		#1		read = 32'd3115648789;
		#1		read = 32'd3134768636;
		#1		read = 32'd3153789755;
		#1		read = 32'd3172710244;
		#1		read = 32'd3191528211;
		#1		read = 32'd3210241775;
		#1		read = 32'd3228849064;
		#1		read = 32'd3247348217;
		#1		read = 32'd3265737385;
		#1		read = 32'd3284014728;
		#1		read = 32'd3302178419;
		#1		read = 32'd3320226642;
		#1		read = 32'd3338157591;
		#1		read = 32'd3355969474;
		#1		read = 32'd3373660509;
		#1		read = 32'd3391228928;
		#1		read = 32'd3408672973;
		#1		read = 32'd3425990900;
		#1		read = 32'd3443180978;
		#1		read = 32'd3460241487;
		#1		read = 32'd3477170721;
		#1		read = 32'd3493966987;
		#1		read = 32'd3510628607;
		#1		read = 32'd3527153913;
		#1		read = 32'd3543541253;
		#1		read = 32'd3559788989;
		#1		read = 32'd3575895495;
		#1		read = 32'd3591859161;
		#1		read = 32'd3607678391;
		#1		read = 32'd3623351603;
		#1		read = 32'd3638877229;
		#1		read = 32'd3654253717;
		#1		read = 32'd3669479529;
		#1		read = 32'd3684553143;
		#1		read = 32'd3699473051;
		#1		read = 32'd3714237762;
		#1		read = 32'd3728845798;
		#1		read = 32'd3743295700;
		#1		read = 32'd3757586021;
		#1		read = 32'd3771715334;
		#1		read = 32'd3785682225;
		#1		read = 32'd3799485297;
		#1		read = 32'd3813123171;
		#1		read = 32'd3826594482;
		#1		read = 32'd3839897884;
		#1		read = 32'd3853032045;
		#1		read = 32'd3865995653;
		#1		read = 32'd3878787411;
		#1		read = 32'd3891406041;
		#1		read = 32'd3903850279;
		#1		read = 32'd3916118883;
		#1		read = 32'd3928210624;
		#1		read = 32'd3940124294;
		#1		read = 32'd3951858701;
		#1		read = 32'd3963412673;
		#1		read = 32'd3974785053;
		#1		read = 32'd3985974704;
		#1		read = 32'd3996980508;
		#1		read = 32'd4007801364;
		#1		read = 32'd4018436190;
		#1		read = 32'd4028883922;
		#1		read = 32'd4039143515;
		#1		read = 32'd4049213944;
		#1		read = 32'd4059094201;
		#1		read = 32'd4068783299;
		#1		read = 32'd4078280269;
		#1		read = 32'd4087584161;
		#1		read = 32'd4096694044;
		#1		read = 32'd4105609008;
		#1		read = 32'd4114328161;
		#1		read = 32'd4122850631;
		#1		read = 32'd4131175566;
		#1		read = 32'd4139302133;
		#1		read = 32'd4147229521;
		#1		read = 32'd4154956935;
		#1		read = 32'd4162483604;
		#1		read = 32'd4169808774;
		#1		read = 32'd4176931714;
		#1		read = 32'd4183851710;
		#1		read = 32'd4190568072;
		#1		read = 32'd4197080126;
		#1		read = 32'd4203387223;
		#1		read = 32'd4209488731;
		#1		read = 32'd4215384040;
		#1		read = 32'd4221072561;
		#1		read = 32'd4226553725;
		#1		read = 32'd4231826983;
		#1		read = 32'd4236891809;
		#1		read = 32'd4241747696;
		#1		read = 32'd4246394158;
		#1		read = 32'd4250830731;
		#1		read = 32'd4255056971;
		#1		read = 32'd4259072455;
		#1		read = 32'd4262876783;
		#1		read = 32'd4266469572;
		#1		read = 32'd4269850465;
		#1		read = 32'd4273019123;
		#1		read = 32'd4275975229;
		#1		read = 32'd4278718488;
		#1		read = 32'd4281248625;
		#1		read = 32'd4283565387;
		#1		read = 32'd4285668543;
		#1		read = 32'd4287557882;
		#1		read = 32'd4289233216;
		#1		read = 32'd4290694376;
		#1		read = 32'd4291941218;
		#1		read = 32'd4292973615;
		#1		read = 32'd4293791465;
		#1		read = 32'd4294394686;
		#1		read = 32'd4294783217;
		#1		read = 32'd4294957021;
		#1		read = 32'd4294916079;
		#1		read = 32'd4294660395;
		#1		read = 32'd4294189996;
		#1		read = 32'd4293504927;
		#1		read = 32'd4292605259;
		#1		read = 32'd4291491080;
		#1		read = 32'd4290162502;
		#1		read = 32'd4288619658;
		#1		read = 32'd4286862702;
		#1		read = 32'd4284891810;
		#1		read = 32'd4282707179;
		#1		read = 32'd4280309028;
		#1		read = 32'd4277697595;
		#1		read = 32'd4274873143;
		#1		read = 32'd4271835954;
		#1		read = 32'd4268586332;
		#1		read = 32'd4265124600;
		#1		read = 32'd4261451107;
		#1		read = 32'd4257566219;
		#1		read = 32'd4253470324;
		#1		read = 32'd4249163832;
		#1		read = 32'd4244647174;
		#1		read = 32'd4239920801;
		#1		read = 32'd4234985186;
		#1		read = 32'd4229840823;
		#1		read = 32'd4224488226;
		#1		read = 32'd4218927931;
		#1		read = 32'd4213160492;
		#1		read = 32'd4207186488;
		#1		read = 32'd4201006515;
		#1		read = 32'd4194621191;
		#1		read = 32'd4188031155;
		#1		read = 32'd4181237067;
		#1		read = 32'd4174239604;
		#1		read = 32'd4167039468;
		#1		read = 32'd4159637378;
		#1		read = 32'd4152034074;
		#1		read = 32'd4144230317;
		#1		read = 32'd4136226887;
		#1		read = 32'd4128024584;
		#1		read = 32'd4119624228;
		#1		read = 32'd4111026661;
		#1		read = 32'd4102232740;
		#1		read = 32'd4093243347;
		#1		read = 32'd4084059379;
		#1		read = 32'd4074681755;
		#1		read = 32'd4065111412;
		#1		read = 32'd4055349309;
		#1		read = 32'd4045396421;
		#1		read = 32'd4035253743;
		#1		read = 32'd4024922289;
		#1		read = 32'd4014403093;
		#1		read = 32'd4003697207;
		#1		read = 32'd3992805701;
		#1		read = 32'd3981729664;
		#1		read = 32'd3970470205;
		#1		read = 32'd3959028448;
		#1		read = 32'd3947405538;
		#1		read = 32'd3935602638;
		#1		read = 32'd3923620927;
		#1		read = 32'd3911461603;
		#1		read = 32'd3899125884;
		#1		read = 32'd3886615002;
		#1		read = 32'd3873930208;
		#1		read = 32'd3861072771;
		#1		read = 32'd3848043976;
		#1		read = 32'd3834845127;
		#1		read = 32'd3821477543;
		#1		read = 32'd3807942561;
		#1		read = 32'd3794241534;
		#1		read = 32'd3780375833;
		#1		read = 32'd3766346844;
		#1		read = 32'd3752155971;
		#1		read = 32'd3737804631;
		#1		read = 32'd3723294261;
		#1		read = 32'd3708626310;
		#1		read = 32'd3693802247;
		#1		read = 32'd3678823554;
		#1		read = 32'd3663691727;
		#1		read = 32'd3648408281;
		#1		read = 32'd3632974744;
		#1		read = 32'd3617392659;
		#1		read = 32'd3601663584;
		#1		read = 32'd3585789093;
		#1		read = 32'd3569770772;
		#1		read = 32'd3553610223;
		#1		read = 32'd3537309064;
		#1		read = 32'd3520868922;
		#1		read = 32'd3504291444;
		#1		read = 32'd3487578285;
		#1		read = 32'd3470731119;
		#1		read = 32'd3453751628;
		#1		read = 32'd3436641512;
		#1		read = 32'd3419402482;
		#1		read = 32'd3402036260;
		#1		read = 32'd3384544585;
		#1		read = 32'd3366929204;
		#1		read = 32'd3349191879;
		#1		read = 32'd3331334385;
		#1		read = 32'd3313358507;
		#1		read = 32'd3295266042;
		#1		read = 32'd3277058800;
		#1		read = 32'd3258738602;
		#1		read = 32'd3240307278;
		#1		read = 32'd3221766674;
		#1		read = 32'd3203118642;
		#1		read = 32'd3184365047;
		#1		read = 32'd3165507765;
		#1		read = 32'd3146548682;
		#1		read = 32'd3127489692;
		#1		read = 32'd3108332703;
		#1		read = 32'd3089079630;
		#1		read = 32'd3069732398;
		#1		read = 32'd3050292942;
		#1		read = 32'd3030763206;
		#1		read = 32'd3011145143;
		#1		read = 32'd2991440714;
		#1		read = 32'd2971651890;
		#1		read = 32'd2951780650;
		#1		read = 32'd2931828981;
		#1		read = 32'd2911798878;
		#1		read = 32'd2891692345;
		#1		read = 32'd2871511391;
		#1		read = 32'd2851258034;
		#1		read = 32'd2830934301;
		#1		read = 32'd2810542224;
		#1		read = 32'd2790083841;
		#1		read = 32'd2769561199;
		#1		read = 32'd2748976349;
		#1		read = 32'd2728331351;
		#1		read = 32'd2707628268;
		#1		read = 32'd2686869172;
		#1		read = 32'd2666056137;
		#1		read = 32'd2645191246;
		#1		read = 32'd2624276584;
		#1		read = 32'd2603314243;
		#1		read = 32'd2582306319;
		#1		read = 32'd2561254914;
		#1		read = 32'd2540162132;
		#1		read = 32'd2519030082;
		#1		read = 32'd2497860878;
		#1		read = 32'd2476656637;
		#1		read = 32'd2455419479;
		#1		read = 32'd2434151527;
		#1		read = 32'd2412854908;
		#1		read = 32'd2391531753;
		#1		read = 32'd2370184193;
		#1		read = 32'd2348814364;
		#1		read = 32'd2327424401;
		#1		read = 32'd2306016445;
		#1		read = 32'd2284592635;
		#1		read = 32'd2263155114;
		#1		read = 32'd2241706027;
		#1		read = 32'd2220247517;
		#1		read = 32'd2198781731;
		#1		read = 32'd2177310816;
		#1		read = 32'd2155836917;
		#1		read = 32'd2134362183;
		#1		read = 32'd2112888762;
		#1		read = 32'd2091418800;
		#1		read = 32'd2069954444;
		#1		read = 32'd2048497841;
		#1		read = 32'd2027051137;
		#1		read = 32'd2005616475;
		#1		read = 32'd1984196001;
		#1		read = 32'd1962791855;
		#1		read = 32'd1941406178;
		#1		read = 32'd1920041108;
		#1		read = 32'd1898698783;
		#1		read = 32'd1877381336;
		#1		read = 32'd1856090899;
		#1		read = 32'd1834829601;
		#1		read = 32'd1813599568;
		#1		read = 32'd1792402923;
		#1		read = 32'd1771241786;
		#1		read = 32'd1750118273;
		#1		read = 32'd1729034496;
		#1		read = 32'd1707992564;
		#1		read = 32'd1686994580;
		#1		read = 32'd1666042645;
		#1		read = 32'd1645138854;
		#1		read = 32'd1624285297;
		#1		read = 32'd1603484059;
		#1		read = 32'd1582737220;
		#1		read = 32'd1562046856;
		#1		read = 32'd1541415035;
		#1		read = 32'd1520843820;
		#1		read = 32'd1500335269;
		#1		read = 32'd1479891432;
		#1		read = 32'd1459514354;
		#1		read = 32'd1439206072;
		#1		read = 32'd1418968617;
		#1		read = 32'd1398804014;
		#1		read = 32'd1378714277;
		#1		read = 32'd1358701417;
		#1		read = 32'd1338767434;
		#1		read = 32'd1318914323;
		#1		read = 32'd1299144067;
		#1		read = 32'd1279458645;
		#1		read = 32'd1259860025;
		#1		read = 32'd1240350166;
		#1		read = 32'd1220931020;
		#1		read = 32'd1201604528;
		#1		read = 32'd1182372623;
		#1		read = 32'd1163237229;
		#1		read = 32'd1144200259;
		#1		read = 32'd1125263616;
		#1		read = 32'd1106429194;
		#1		read = 32'd1087698877;
		#1		read = 32'd1069074537;
		#1		read = 32'd1050558037;
		#1		read = 32'd1032151229;
		#1		read = 32'd1013855954;
		#1		read = 32'd995674040;
		#1		read = 32'd977607306;
		#1		read = 32'd959657559;
		#1		read = 32'd941826593;
		#1		read = 32'd924116192;
		#1		read = 32'd906528127;
		#1		read = 32'd889064157;
		#1		read = 32'd871726027;
		#1		read = 32'd854515472;
		#1		read = 32'd837434213;
		#1		read = 32'd820483957;
		#1		read = 32'd803666401;
		#1		read = 32'd786983225;
		#1		read = 32'd770436098;
		#1		read = 32'd754026674;
		#1		read = 32'd737756595;
		#1		read = 32'd721627488;
		#1		read = 32'd705640965;
		#1		read = 32'd689798625;
		#1		read = 32'd674102053;
		#1		read = 32'd658552817;
		#1		read = 32'd643152473;
		#1		read = 32'd627902561;
		#1		read = 32'd612804606;
		#1		read = 32'd597860118;
		#1		read = 32'd583070590;
		#1		read = 32'd568437503;
		#1		read = 32'd553962319;
		#1		read = 32'd539646485;
		#1		read = 32'd525491434;
		#1		read = 32'd511498581;
		#1		read = 32'd497669325;
		#1		read = 32'd484005049;
		#1		read = 32'd470507120;
		#1		read = 32'd457176887;
		#1		read = 32'd444015683;
		#1		read = 32'd431024825;
		#1		read = 32'd418205610;
		#1		read = 32'd405559323;
		#1		read = 32'd393087226;
		#1		read = 32'd380790568;
		#1		read = 32'd368670577;
		#1		read = 32'd356728466;
		#1		read = 32'd344965429;
		#1		read = 32'd333382643;
		#1		read = 32'd321981265;
		#1		read = 32'd310762436;
		#1		read = 32'd299727277;
		#1		read = 32'd288876892;
		#1		read = 32'd278212367;
		#1		read = 32'd267734767;
		#1		read = 32'd257445141;
		#1		read = 32'd247344516;
		#1		read = 32'd237433905;
		#1		read = 32'd227714296;
		#1		read = 32'd218186663;
		#1		read = 32'd208851958;
		#1		read = 32'd199711114;
		#1		read = 32'd190765046;
		#1		read = 32'd182014649;
		#1		read = 32'd173460796;
		#1		read = 32'd165104345;
		#1		read = 32'd156946129;
		#1		read = 32'd148986966;
		#1		read = 32'd141227650;
		#1		read = 32'd133668959;
		#1		read = 32'd126311647;
		#1		read = 32'd119156451;
		#1		read = 32'd112204086;
		#1		read = 32'd105455247;
		#1		read = 32'd98910609;
		#1		read = 32'd92570827;
		#1		read = 32'd86436534;
		#1		read = 32'd80508345;
		#1		read = 32'd74786851;
		#1		read = 32'd69272625;
		#1		read = 32'd63966219;
		#1		read = 32'd58868162;
		#1		read = 32'd53978966;
		#1		read = 32'd49299118;
		#1		read = 32'd44829087;
		#1		read = 32'd40569319;
		#1		read = 32'd36520241;
		#1		read = 32'd32682258;
		#1		read = 32'd29055753;
		#1		read = 32'd25641089;
		#1		read = 32'd22438608;
		#1		read = 32'd19448629;
		#1		read = 32'd16671453;
		#1		read = 32'd14107355;
		#1		read = 32'd11756594;
		#1		read = 32'd9619403;
		#1		read = 32'd7695997;
		#1		read = 32'd5986568;
		#1		read = 32'd4491287;
		#1		read = 32'd3210303;
		#1		read = 32'd2143745;
		#1		read = 32'd1291719;
		#1		read = 32'd654310;
		#1		read = 32'd231583;
		#1		read = 32'd23579;
		#1		read = 32'd30319;
		#1		read = 32'd251803;
		#1		read = 32'd688008;
		#1		read = 32'd1338891;
		#1		read = 32'd2204387;
		#1		read = 32'd3284409;
		#1		read = 32'd4578849;
		#1		read = 32'd6087577;
		#1		read = 32'd7810444;
		#1		read = 32'd9747276;
		#1		read = 32'd11897880;
		#1		read = 32'd14262040;
		#1		read = 32'd16839521;
		#1		read = 32'd19630065;
		#1		read = 32'd22633392;
		#1		read = 32'd25849203;
		#1		read = 32'd29277175;
		#1		read = 32'd32916966;
		#1		read = 32'd36768212;
		#1		read = 32'd40830528;
		#1		read = 32'd45103507;
		#1		read = 32'd49586723;
		#1		read = 32'd54279726;
		#1		read = 32'd59182048;
		#1		read = 32'd64293199;
		#1		read = 32'd69612667;
		#1		read = 32'd75139920;
		#1		read = 32'd80874406;
		#1		read = 32'd86815551;
		#1		read = 32'd92962761;
		#1		read = 32'd99315422;
		#1		read = 32'd105872898;
		#1		read = 32'd112634533;
		#1		read = 32'd119599651;
		#1		read = 32'd126767556;
		#1		read = 32'd134137531;
		#1		read = 32'd141708839;
		#1		read = 32'd149480722;
		#1		read = 32'd157452405;
		#1		read = 32'd165623088;
		#1		read = 32'd173991957;
		#1		read = 32'd182558172;
		#1		read = 32'd191320879;
		#1		read = 32'd200279200;
		#1		read = 32'd209432240;
		#1		read = 32'd218779084;
		#1		read = 32'd228318796;
		#1		read = 32'd238050424;
		#1		read = 32'd247972993;
		#1		read = 32'd258085511;
		#1		read = 32'd268386968;
		#1		read = 32'd278876333;
		#1		read = 32'd289552557;
		#1		read = 32'd300414573;
		#1		read = 32'd311461294;
		#1		read = 32'd322691615;
		#1		read = 32'd334104415;
		#1		read = 32'd345698550;
		#1		read = 32'd357472863;
		#1		read = 32'd369426176;
		#1		read = 32'd381557292;
		#1		read = 32'd393865000;
		#1		read = 32'd406348068;
		#1		read = 32'd419005249;
		#1		read = 32'd431835275;
		#1		read = 32'd444836865;
		#1		read = 32'd458008719;
		#1		read = 32'd471349518;
		#1		read = 32'd484857930;
		#1		read = 32'd498532602;
		#1		read = 32'd512372169;
		#1		read = 32'd526375245;
		#1		read = 32'd540540431;
		#1		read = 32'd554866309;
		#1		read = 32'd569351448;
		#1		read = 32'd583994399;
		#1		read = 32'd598793698;
		#1		read = 32'd613747864;
		#1		read = 32'd628855403;
		#1		read = 32'd644114803;
		#1		read = 32'd659524539;
		#1		read = 32'd675083069;
		#1		read = 32'd690788839;
		#1		read = 32'd706640276;
		#1		read = 32'd722635797;
		#1		read = 32'd738773801;
		#1		read = 32'd755052675;
		#1		read = 32'd771470791;
		#1		read = 32'd788026507;
		#1		read = 32'd804718168;
		#1		read = 32'd821544104;
		#1		read = 32'd838502633;
		#1		read = 32'd855592060;
		#1		read = 32'd872810674;
		#1		read = 32'd890156754;
		#1		read = 32'd907628566;
		#1		read = 32'd925224363;
		#1		read = 32'd942942384;
		#1		read = 32'd960780858;
		#1		read = 32'd978738002;
		#1		read = 32'd996812020;
		#1		read = 32'd1015001103;
		#1		read = 32'd1033303434;
		#1		read = 32'd1051717182;
		#1		read = 32'd1070240506;
		#1		read = 32'd1088871553;
		#1		read = 32'd1107608461;
		#1		read = 32'd1126449355;
		#1		read = 32'd1145392351;
		#1		read = 32'd1164435556;
		#1		read = 32'd1183577065;
		#1		read = 32'd1202814964;
		#1		read = 32'd1222147329;
		#1		read = 32'd1241572227;
		#1		read = 32'd1261087715;
		#1		read = 32'd1280691842;
		#1		read = 32'd1300382648;
		#1		read = 32'd1320158163;
		#1		read = 32'd1340016409;
		#1		read = 32'd1359955402;
		#1		read = 32'd1379973147;
		#1		read = 32'd1400067642;
		#1		read = 32'd1420236879;
		#1		read = 32'd1440478839;
		#1		read = 32'd1460791500;
		#1		read = 32'd1481172829;
		#1		read = 32'd1501620788;
		#1		read = 32'd1522133333;
		#1		read = 32'd1542708413;
		#1		read = 32'd1563343970;
		#1		read = 32'd1584037940;
		#1		read = 32'd1604788254;
		#1		read = 32'd1625592838;
		#1		read = 32'd1646449610;
		#1		read = 32'd1667356485;
		#1		read = 32'd1688311372;
		#1		read = 32'd1709312177;
		#1		read = 32'd1730356798;
		#1		read = 32'd1751443131;
		#1		read = 32'd1772569068;
		#1		read = 32'd1793732496;
		#1		read = 32'd1814931299;
		#1		read = 32'd1836163357;
		#1		read = 32'd1857426547;
		#1		read = 32'd1878718742;
		#1		read = 32'd1900037814;
		#1		read = 32'd1921381630;
		#1		read = 32'd1942748056;
		#1		read = 32'd1964134955;
		#1		read = 32'd1985540189;
		#1		read = 32'd2006961617;
		#1		read = 32'd2028397097;
		#1		read = 32'd2049844486;
		#1		read = 32'd2071301639;
		#1		read = 32'd2092766410;
		#1		read = 32'd2114236652;
		#1		read = 32'd2135710219;
		#1		read = 32'd2157184964;
		#1		read = 32'd2178658738;
		#1		read = 32'd2200129395;
		#1		read = 32'd2221594787;
		#1		read = 32'd2243052769;
		#1		read = 32'd2264501193;
		#1		read = 32'd2285937916;
		#1		read = 32'd2307360794;
		#1		read = 32'd2328767683;
		#1		read = 32'd2350156445;
		#1		read = 32'd2371524940;
		#1		read = 32'd2392871030;
		#1		read = 32'd2414192582;
		#1		read = 32'd2435487464;
		#1		read = 32'd2456753545;
		#1		read = 32'd2477988700;
		#1		read = 32'd2499190804;
		#1		read = 32'd2520357738;
		#1		read = 32'd2541487385;
		#1		read = 32'd2562577631;
		#1		read = 32'd2583626369;
		#1		read = 32'd2604631493;
		#1		read = 32'd2625590902;
		#1		read = 32'd2646502501;
		#1		read = 32'd2667364199;
		#1		read = 32'd2688173909;
		#1		read = 32'd2708929550;
		#1		read = 32'd2729629048;
		#1		read = 32'd2750270331;
		#1		read = 32'd2770851336;
		#1		read = 32'd2791370005;
		#1		read = 32'd2811824285;
		#1		read = 32'd2832212133;
		#1		read = 32'd2852531507;
		#1		read = 32'd2872780378;
		#1		read = 32'd2892956720;
		#1		read = 32'd2913058515;
		#1		read = 32'd2933083753;
		#1		read = 32'd2953030432;
		#1		read = 32'd2972896556;
		#1		read = 32'd2992680141;
		#1		read = 32'd3012379206;
		#1		read = 32'd3031991782;
		#1		read = 32'd3051515908;
		#1		read = 32'd3070949632;
		#1		read = 32'd3090291010;
		#1		read = 32'd3109538108;
		#1		read = 32'd3128689002;
		#1		read = 32'd3147741775;
		#1		read = 32'd3166694524;
		#1		read = 32'd3185545352;
		#1		read = 32'd3204292376;
		#1		read = 32'd3222933719;
		#1		read = 32'd3241467518;
		#1		read = 32'd3259891919;
		#1		read = 32'd3278205081;
		#1		read = 32'd3296405172;
		#1		read = 32'd3314490371;
		#1		read = 32'd3332458870;
		#1		read = 32'd3350308873;
		#1		read = 32'd3368038595;
		#1		read = 32'd3385646262;
		#1		read = 32'd3403130114;
		#1		read = 32'd3420488402;
		#1		read = 32'd3437719391;
		#1		read = 32'd3454821357;
		#1		read = 32'd3471792591;
		#1		read = 32'd3488631395;
		#1		read = 32'd3505336085;
		#1		read = 32'd3521904991;
		#1		read = 32'd3538336456;
		#1		read = 32'd3554628837;
		#1		read = 32'd3570780504;
		#1		read = 32'd3586789844;
		#1		read = 32'd3602655253;
		#1		read = 32'd3618375147;
		#1		read = 32'd3633947953;
		#1		read = 32'd3649372113;
		#1		read = 32'd3664646086;
		#1		read = 32'd3679768344;
		#1		read = 32'd3694737375;
		#1		read = 32'd3709551682;
		#1		read = 32'd3724209783;
		#1		read = 32'd3738710213;
		#1		read = 32'd3753051522;
		#1		read = 32'd3767232275;
		#1		read = 32'd3781251055;
		#1		read = 32'd3795106459;
		#1		read = 32'd3808797102;
		#1		read = 32'd3822321616;
		#1		read = 32'd3835678647;
		#1		read = 32'd3848866860;
		#1		read = 32'd3861884936;
		#1		read = 32'd3874731573;
		#1		read = 32'd3887405487;
		#1		read = 32'd3899905410;
		#1		read = 32'd3912230093;
		#1		read = 32'd3924378302;
		#1		read = 32'd3936348824;
		#1		read = 32'd3948140460;
		#1		read = 32'd3959752032;
		#1		read = 32'd3971182379;
		#1		read = 32'd3982430358;
		#1		read = 32'd3993494843;
		#1		read = 32'd4004374729;
		#1		read = 32'd4015068927;
		#1		read = 32'd4025576368;
		#1		read = 32'd4035896002;
		#1		read = 32'd4046026795;
		#1		read = 32'd4055967737;
		#1		read = 32'd4065717831;
		#1		read = 32'd4075276103;
		#1		read = 32'd4084641598;
		#1		read = 32'd4093813379;
		#1		read = 32'd4102790528;
		#1		read = 32'd4111572148;
		#1		read = 32'd4120157361;
		#1		read = 32'd4128545309;
		#1		read = 32'd4136735152;
		#1		read = 32'd4144726071;
		#1		read = 32'd4152517268;
		#1		read = 32'd4160107963;
		#1		read = 32'd4167497397;
		#1		read = 32'd4174684831;
		#1		read = 32'd4181669548;
		#1		read = 32'd4188450847;
		#1		read = 32'd4195028051;
		#1		read = 32'd4201400503;
		#1		read = 32'd4207567564;
		#1		read = 32'd4213528619;
		#1		read = 32'd4219283071;
		#1		read = 32'd4224830345;
		#1		read = 32'd4230169886;
		#1		read = 32'd4235301160;
		#1		read = 32'd4240223654;
		#1		read = 32'd4244936876;
		#1		read = 32'd4249440354;
		#1		read = 32'd4253733638;
		#1		read = 32'd4257816299;
		#1		read = 32'd4261687929;
		#1		read = 32'd4265348140;
		#1		read = 32'd4268796566;
		#1		read = 32'd4272032863;
		#1		read = 32'd4275056706;
		#1		read = 32'd4277867794;
		#1		read = 32'd4280465845;
		#1		read = 32'd4282850600;
		#1		read = 32'd4285021820;
		#1		read = 32'd4286979288;
		#1		read = 32'd4288722808;
		#1		read = 32'd4290252206;
		#1		read = 32'd4291567329;
		#1		read = 32'd4292668046;
		#1		read = 32'd4293554245;
		#1		read = 32'd4294225840;
		#1		read = 32'd4294682762;
		#1		read = 32'd4294924966;
		#1		read = 32'd4294952427;
		#1		read = 32'd4294765144;
		#1		read = 32'd4294363134;
		#1		read = 32'd4293746438;
		#1		read = 32'd4292915117;
		#1		read = 32'd4291869256;
		#1		read = 32'd4290608957;
		#1		read = 32'd4289134347;
		#1		read = 32'd4287445575;
		#1		read = 32'd4285542808;
		#1		read = 32'd4283426236;
		#1		read = 32'd4281096073;
		#1		read = 32'd4278552549;
		#1		read = 32'd4275795921;
		#1		read = 32'd4272826463;
		#1		read = 32'd4269644473;
		#1		read = 32'd4266250269;
		#1		read = 32'd4262644189;
		#1		read = 32'd4258826595;
		#1		read = 32'd4254797869;
		#1		read = 32'd4250558413;
		#1		read = 32'd4246108651;
		#1		read = 32'd4241449029;
		#1		read = 32'd4236580012;
		#1		read = 32'd4231502087;
		#1		read = 32'd4226215761;
		#1		read = 32'd4220721565;
		#1		read = 32'd4215020046;
		#1		read = 32'd4209111775;
		#1		read = 32'd4202997343;
		#1		read = 32'd4196677362;
		#1		read = 32'd4190152463;
		#1		read = 32'd4183423298;
		#1		read = 32'd4176490542;
		#1		read = 32'd4169354886;
		#1		read = 32'd4162017045;
		#1		read = 32'd4154477753;
		#1		read = 32'd4146737762;
		#1		read = 32'd4138797848;
		#1		read = 32'd4130658804;
		#1		read = 32'd4122321444;
		#1		read = 32'd4113786603;
		#1		read = 32'd4105055132;
		#1		read = 32'd4096127906;
		#1		read = 32'd4087005817;
		#1		read = 32'd4077689778;
		#1		read = 32'd4068180719;
		#1		read = 32'd4058479592;
		#1		read = 32'd4048587368;
		#1		read = 32'd4038505034;
		#1		read = 32'd4028233601;
		#1		read = 32'd4017774093;
		#1		read = 32'd4007127558;
		#1		read = 32'd3996295061;
		#1		read = 32'd3985277683;
		#1		read = 32'd3974076528;
		#1		read = 32'd3962692715;
		#1		read = 32'd3951127383;
		#1		read = 32'd3939381688;
		#1		read = 32'd3927456804;
		#1		read = 32'd3915353925;
		#1		read = 32'd3903074260;
		#1		read = 32'd3890619037;
		#1		read = 32'd3877989503;
		#1		read = 32'd3865186919;
		#1		read = 32'd3852212566;
		#1		read = 32'd3839067742;
		#1		read = 32'd3825753761;
		#1		read = 32'd3812271955;
		#1		read = 32'd3798623670;
		#1		read = 32'd3784810274;
		#1		read = 32'd3770833146;
		#1		read = 32'd3756693684;
		#1		read = 32'd3742393303;
		#1		read = 32'd3727933432;
		#1		read = 32'd3713315517;
		#1		read = 32'd3698541020;
		#1		read = 32'd3683611420;
		#1		read = 32'd3668528207;
		#1		read = 32'd3653292891;
		#1		read = 32'd3637906996;
		#1		read = 32'd3622372060;
		#1		read = 32'd3606689636;
		#1		read = 32'd3590861292;
		#1		read = 32'd3574888612;
		#1		read = 32'd3558773193;
		#1		read = 32'd3542516646;
		#1		read = 32'd3526120597;
		#1		read = 32'd3509586685;
		#1		read = 32'd3492916564;
		#1		read = 32'd3476111901;
		#1		read = 32'd3459174376;
		#1		read = 32'd3442105684;
		#1		read = 32'd3424907530;
		#1		read = 32'd3407581634;
		#1		read = 32'd3390129730;
		#1		read = 32'd3372553563;
		#1		read = 32'd3354854889;
		#1		read = 32'd3337035480;
		#1		read = 32'd3319097116;
		#1		read = 32'd3301041592;
		#1		read = 32'd3282870713;
		#1		read = 32'd3264586296;
		#1		read = 32'd3246190170;
		#1		read = 32'd3227684174;
		#1		read = 32'd3209070159;
		#1		read = 32'd3190349986;
		#1		read = 32'd3171525528;
		#1		read = 32'd3152598666;
		#1		read = 32'd3133571293;
		#1		read = 32'd3114445313;
		#1		read = 32'd3095222637;
		#1		read = 32'd3075905188;
		#1		read = 32'd3056494898;
		#1		read = 32'd3036993707;
		#1		read = 32'd3017403566;
		#1		read = 32'd2997726434;
		#1		read = 32'd2977964278;
		#1		read = 32'd2958119075;
		#1		read = 32'd2938192809;
		#1		read = 32'd2918187473;
		#1		read = 32'd2898105067;
		#1		read = 32'd2877947599;
		#1		read = 32'd2857717086;
		#1		read = 32'd2837415550;
		#1		read = 32'd2817045021;
		#1		read = 32'd2796607537;
		#1		read = 32'd2776105140;
		#1		read = 32'd2755539883;
		#1		read = 32'd2734913820;
		#1		read = 32'd2714229014;
		#1		read = 32'd2693487535;
		#1		read = 32'd2672691456;
		#1		read = 32'd2651842856;
		#1		read = 32'd2630943821;
		#1		read = 32'd2609996440;
		#1		read = 32'd2589002808;
		#1		read = 32'd2567965025;
		#1		read = 32'd2546885194;
		#1		read = 32'd2525765423;
		#1		read = 32'd2504607824;
		#1		read = 32'd2483414513;
		#1		read = 32'd2462187609;
		#1		read = 32'd2440929236;
		#1		read = 32'd2419641517;
		#1		read = 32'd2398326584;
		#1		read = 32'd2376986566;
		#1		read = 32'd2355623598;
		#1		read = 32'd2334239816;
		#1		read = 32'd2312837359;
		#1		read = 32'd2291418367;
		#1		read = 32'd2269984981;
		#1		read = 32'd2248539345;
		#1		read = 32'd2227083604;
		#1		read = 32'd2205619903;
		#1		read = 32'd2184150388;
		#1		read = 32'd2162677206;
		#1		read = 32'd2141202506;
		#1		read = 32'd2119728433;
		#1		read = 32'd2098257136;
		#1		read = 32'd2076790761;
		#1		read = 32'd2055331456;
		#1		read = 32'd2033881366;
		#1		read = 32'd2012442636;
		#1		read = 32'd1991017410;
		#1		read = 32'd1969607830;
		#1		read = 32'd1948216038;
		#1		read = 32'd1926844173;
		#1		read = 32'd1905494371;
		#1		read = 32'd1884168768;
		#1		read = 32'd1862869496;
		#1		read = 32'd1841598685;
		#1		read = 32'd1820358463;
		#1		read = 32'd1799150953;
		#1		read = 32'd1777978276;
		#1		read = 32'd1756842549;
		#1		read = 32'd1735745886;
		#1		read = 32'd1714690396;
		#1		read = 32'd1693678185;
		#1		read = 32'd1672711355;
		#1		read = 32'd1651792001;
		#1		read = 32'd1630922216;
		#1		read = 32'd1610104087;
		#1		read = 32'd1589339695;
		#1		read = 32'd1568631117;
		#1		read = 32'd1547980424;
		#1		read = 32'd1527389681;
		#1		read = 32'd1506860947;
		#1		read = 32'd1486396274;
		#1		read = 32'd1465997710;
		#1		read = 32'd1445667293;
		#1		read = 32'd1425407058;
		#1		read = 32'd1405219030;
		#1		read = 32'd1385105227;
		#1		read = 32'd1365067662;
		#1		read = 32'd1345108338;
		#1		read = 32'd1325229250;
		#1		read = 32'd1305432388;
		#1		read = 32'd1285719729;
		#1		read = 32'd1266093247;
		#1		read = 32'd1246554903;
		#1		read = 32'd1227106650;
		#1		read = 32'd1207750435;
		#1		read = 32'd1188488193;
		#1		read = 32'd1169321849;
		#1		read = 32'd1150253320;
		#1		read = 32'd1131284514;
		#1		read = 32'd1112417326;
		#1		read = 32'd1093653645;
		#1		read = 32'd1074995345;
		#1		read = 32'd1056444294;
		#1		read = 32'd1038002346;
		#1		read = 32'd1019671344;
		#1		read = 32'd1001453123;
		#1		read = 32'd983349505;
		#1		read = 32'd965362298;
		#1		read = 32'd947493303;
		#1		read = 32'd929744306;
		#1		read = 32'd912117081;
		#1		read = 32'd894613393;
		#1		read = 32'd877234990;
		#1		read = 32'd859983611;
		#1		read = 32'd842860981;
		#1		read = 32'd825868812;
		#1		read = 32'd809008804;
		#1		read = 32'd792282642;
		#1		read = 32'd775691999;
		#1		read = 32'd759238534;
		#1		read = 32'd742923892;
		#1		read = 32'd726749705;
		#1		read = 32'd710717591;
		#1		read = 32'd694829152;
		#1		read = 32'd679085977;
		#1		read = 32'd663489640;
		#1		read = 32'd648041702;
		#1		read = 32'd632743706;
		#1		read = 32'd617597184;
		#1		read = 32'd602603649;
		#1		read = 32'd587764600;
		#1		read = 32'd573081522;
		#1		read = 32'd558555883;
		#1		read = 32'd544189135;
		#1		read = 32'd529982716;
		#1		read = 32'd515938045;
		#1		read = 32'd502056528;
		#1		read = 32'd488339552;
		#1		read = 32'd474788488;
		#1		read = 32'd461404693;
		#1		read = 32'd448189505;
		#1		read = 32'd435144244;
		#1		read = 32'd422270216;
		#1		read = 32'd409568708;
		#1		read = 32'd397040990;
		#1		read = 32'd384688315;
		#1		read = 32'd372511918;
		#1		read = 32'd360513016;
		#1		read = 32'd348692810;
		#1		read = 32'd337052482;
		#1		read = 32'd325593195;
		#1		read = 32'd314316096;
		#1		read = 32'd303222312;
		#1		read = 32'd292312952;
		#1		read = 32'd281589109;
		#1		read = 32'd271051853;
		#1		read = 32'd260702238;
		#1		read = 32'd250541300;
		#1		read = 32'd240570055;
		#1		read = 32'd230789500;
		#1		read = 32'd221200612;
		#1		read = 32'd211804352;
		#1		read = 32'd202601657;
		#1		read = 32'd193593449;
		#1		read = 32'd184780629;
		#1		read = 32'd176164077;
		#1		read = 32'd167744655;
		#1		read = 32'd159523206;
		#1		read = 32'd151500551;
		#1		read = 32'd143677493;
		#1		read = 32'd136054813;
		#1		read = 32'd128633275;
		#1		read = 32'd121413620;
		#1		read = 32'd114396571;
		#1		read = 32'd107582828;
		#1		read = 32'd100973074;
		#1		read = 32'd94567970;
		#1		read = 32'd88368155;
		#1		read = 32'd82374250;
		#1		read = 32'd76586854;
		#1		read = 32'd71006546;
		#1		read = 32'd65633884;
		#1		read = 32'd60469405;
		#1		read = 32'd55513626;
		#1		read = 32'd50767043;
		#1		read = 32'd46230129;
		#1		read = 32'd41903339;
		#1		read = 32'd37787105;
		#1		read = 32'd33881839;
		#1		read = 32'd30187931;
		#1		read = 32'd26705752;
		#1		read = 32'd23435648;
		#1		read = 32'd20377947;
		#1		read = 32'd17532955;
		#1		read = 32'd14900956;
		#1		read = 32'd12482214;
		#1		read = 32'd10276971;
		#1		read = 32'd8285446;
		#1		read = 32'd6507839;
		#1		read = 32'd4944328;
		#1		read = 32'd3595069;
		#1		read = 32'd2460197;
		#1		read = 32'd1539826;
		#1		read = 32'd834047;
		#1		read = 32'd342931;
		#1		read = 32'd66528;
		#1		read = 32'd4865;
		#1		read = 32'd157948;
		#1		read = 32'd525761;
		#1		read = 32'd1108269;
		#1		read = 32'd1905412;
		#1		read = 32'd2917111;
		#1		read = 32'd4143266;
		#1		read = 32'd5583752;
		#1		read = 32'd7238427;
		#1		read = 32'd9107124;
		#1		read = 32'd11189657;
		#1		read = 32'd13485818;
		#1		read = 32'd15995377;
		#1		read = 32'd18718083;
		#1		read = 32'd21653664;
		#1		read = 32'd24801826;
		#1		read = 32'd28162254;
		#1		read = 32'd31734613;
		#1		read = 32'd35518545;
		#1		read = 32'd39513671;
		#1		read = 32'd43719593;
		#1		read = 32'd48135890;
		#1		read = 32'd52762119;
		#1		read = 32'd57597819;
		#1		read = 32'd62642506;
		#1		read = 32'd67895675;
		#1		read = 32'd73356802;
		#1		read = 32'd79025339;
		#1		read = 32'd84900720;
		#1		read = 32'd90982358;
		#1		read = 32'd97269644;
		#1		read = 32'd103761950;
		#1		read = 32'd110458627;
		#1		read = 32'd117359004;
		#1		read = 32'd124462392;
		#1		read = 32'd131768080;
		#1		read = 32'd139275339;
		#1		read = 32'd146983416;
		#1		read = 32'd154891542;
		#1		read = 32'd162998926;
		#1		read = 32'd171304756;
		#1		read = 32'd179808202;
		#1		read = 32'd188508415;
		#1		read = 32'd197404523;
		#1		read = 32'd206495637;
		#1		read = 32'd215780849;
		#1		read = 32'd225259230;
		#1		read = 32'd234929831;
		#1		read = 32'd244791686;
		#1		read = 32'd254843808;
		#1		read = 32'd265085194;
		#1		read = 32'd275514817;
		#1		read = 32'd286131636;
		#1		read = 32'd296934588;
		#1		read = 32'd307922593;
		#1		read = 32'd319094554;
		#1		read = 32'd330449351;
		#1		read = 32'd341985851;
		#1		read = 32'd353702899;
		#1		read = 32'd365599323;
		#1		read = 32'd377673934;
		#1		read = 32'd389925525;
		#1		read = 32'd402352870;
		#1		read = 32'd414954727;
		#1		read = 32'd427729836;
		#1		read = 32'd440676918;
		#1		read = 32'd453794679;
		#1		read = 32'd467081808;
		#1		read = 32'd480536976;
		#1		read = 32'd494158837;
		#1		read = 32'd507946029;
		#1		read = 32'd521897174;
		#1		read = 32'd536010875;
		#1		read = 32'd550285723;
		#1		read = 32'd564720289;
		#1		read = 32'd579313130;
		#1		read = 32'd594062787;
		#1		read = 32'd608967785;
		#1		read = 32'd624026633;
		#1		read = 32'd639237826;
		#1		read = 32'd654599841;
		#1		read = 32'd670111144;
		#1		read = 32'd685770183;
		#1		read = 32'd701575392;
		#1		read = 32'd717525191;
		#1		read = 32'd733617985;
		#1		read = 32'd749852163;
		#1		read = 32'd766226104;
		#1		read = 32'd782738169;
		#1		read = 32'd799386708;
		#1		read = 32'd816170055;
		#1		read = 32'd833086533;
		#1		read = 32'd850134449;
		#1		read = 32'd867312099;
		#1		read = 32'd884617765;
		#1		read = 32'd902049717;
		#1		read = 32'd919606211;
		#1		read = 32'd937285492;
		#1		read = 32'd955085791;
		#1		read = 32'd973005330;
		#1		read = 32'd991042315;
		#1		read = 32'd1009194943;
		#1		read = 32'd1027461399;
		#1		read = 32'd1045839857;
		#1		read = 32'd1064328478;
		#1		read = 32'd1082925414;
		#1		read = 32'd1101628804;
		#1		read = 32'd1120436779;
		#1		read = 32'd1139347458;
		#1		read = 32'd1158358950;
		#1		read = 32'd1177469354;
		#1		read = 32'd1196676758;
		#1		read = 32'd1215979242;
		#1		read = 32'd1235374875;
		#1		read = 32'd1254861719;
		#1		read = 32'd1274437824;
		#1		read = 32'd1294101233;
		#1		read = 32'd1313849980;
		#1		read = 32'd1333682089;
		#1		read = 32'd1353595578;
		#1		read = 32'd1373588455;
		#1		read = 32'd1393658720;
		#1		read = 32'd1413804368;
		#1		read = 32'd1434023383;
		#1		read = 32'd1454313743;
		#1		read = 32'd1474673420;
		#1		read = 32'd1495100377;
		#1		read = 32'd1515592572;
		#1		read = 32'd1536147956;
		#1		read = 32'd1556764473;
		#1		read = 32'd1577440061;
		#1		read = 32'd1598172653;
		#1		read = 32'd1618960175;
		#1		read = 32'd1639800550;
		#1		read = 32'd1660691692;
		#1		read = 32'd1681631513;
		#1		read = 32'd1702617919;
		#1		read = 32'd1723648812;
		#1		read = 32'd1744722087;
		#1		read = 32'd1765835638;
		#1		read = 32'd1786987354;
		#1		read = 32'd1808175119;
		#1		read = 32'd1829396814;
		#1		read = 32'd1850650318;
		#1		read = 32'd1871933505;
		#1		read = 32'd1893244247;
		#1		read = 32'd1914580413;
		#1		read = 32'd1935939868;
		#1		read = 32'd1957320478;
		#1		read = 32'd1978720104;
		#1		read = 32'd2000136607;
		#1		read = 32'd2021567844;
		#1		read = 32'd2043011672;
		#1		read = 32'd2064465947;
		#1		read = 32'd2085928524;
		#1		read = 32'd2107397257;
		#1		read = 32'd2128869998;
		#1		read = 32'd2150344601;
		#1		read = 32'd2171818917;
		#1		read = 32'd2193290800;
		#1		read = 32'd2214758103;
		#1		read = 32'd2236218677;
		#1		read = 32'd2257670379;
		#1		read = 32'd2279111062;
		#1		read = 32'd2300538582;
		#1		read = 32'd2321950797;
		#1		read = 32'd2343345565;
		#1		read = 32'd2364720748;
		#1		read = 32'd2386074206;
		#1		read = 32'd2407403806;
		#1		read = 32'd2428707414;
		#1		read = 32'd2449982900;
		#1		read = 32'd2471228137;
		#1		read = 32'd2492440999;
		#1		read = 32'd2513619365;
		#1		read = 32'd2534761119;
		#1		read = 32'd2555864145;
		#1		read = 32'd2576926333;
		#1		read = 32'd2597945577;
		#1		read = 32'd2618919776;
		#1		read = 32'd2639846831;
		#1		read = 32'd2660724650;
		#1		read = 32'd2681551146;
		#1		read = 32'd2702324236;
		#1		read = 32'd2723041841;
		#1		read = 32'd2743701892;
		#1		read = 32'd2764302321;
		#1		read = 32'd2784841069;
		#1		read = 32'd2805316082;
		#1		read = 32'd2825725311;
		#1		read = 32'd2846066718;
		#1		read = 32'd2866338266;
		#1		read = 32'd2886537930;
		#1		read = 32'd2906663689;
		#1		read = 32'd2926713530;
		#1		read = 32'd2946685450;
		#1		read = 32'd2966577449;
		#1		read = 32'd2986387540;
		#1		read = 32'd3006113742;
		#1		read = 32'd3025754081;
		#1		read = 32'd3045306593;
		#1		read = 32'd3064769324;
		#1		read = 32'd3084140328;
		#1		read = 32'd3103417666;
		#1		read = 32'd3122599412;
		#1		read = 32'd3141683647;
		#1		read = 32'd3160668463;
		#1		read = 32'd3179551961;
		#1		read = 32'd3198332254;
		#1		read = 32'd3217007462;
		#1		read = 32'd3235575719;
		#1		read = 32'd3254035167;
		#1		read = 32'd3272383962;
		#1		read = 32'd3290620267;
		#1		read = 32'd3308742259;
		#1		read = 32'd3326748127;
		#1		read = 32'd3344636069;
		#1		read = 32'd3362404297;
		#1		read = 32'd3380051034;
		#1		read = 32'd3397574515;
		#1		read = 32'd3414972988;
		#1		read = 32'd3432244713;
		#1		read = 32'd3449387963;
		#1		read = 32'd3466401024;
		#1		read = 32'd3483282194;
		#1		read = 32'd3500029786;
		#1		read = 32'd3516642124;
		#1		read = 32'd3533117547;
		#1		read = 32'd3549454408;
		#1		read = 32'd3565651073;
		#1		read = 32'd3581705922;
		#1		read = 32'd3597617351;
		#1		read = 32'd3613383767;
		#1		read = 32'd3629003595;
		#1		read = 32'd3644475272;
		#1		read = 32'd3659797251;
		#1		read = 32'd3674967999;
		#1		read = 32'd3689986001;
		#1		read = 32'd3704849754;
		#1		read = 32'd3719557771;
		#1		read = 32'd3734108582;
		#1		read = 32'd3748500732;
		#1		read = 32'd3762732782;
		#1		read = 32'd3776803308;
		#1		read = 32'd3790710904;
		#1		read = 32'd3804454178;
		#1		read = 32'd3818031756;
		#1		read = 32'd3831442281;
		#1		read = 32'd3844684412;
		#1		read = 32'd3857756824;
		#1		read = 32'd3870658210;
		#1		read = 32'd3883387280;
		#1		read = 32'd3895942761;
		#1		read = 32'd3908323398;
		#1		read = 32'd3920527952;
		#1		read = 32'd3932555203;
		#1		read = 32'd3944403949;
		#1		read = 32'd3956073004;
		#1		read = 32'd3967561202;
		#1		read = 32'd3978867393;
		#1		read = 32'd3989990447;
		#1		read = 32'd4000929253;
		#1		read = 32'd4011682715;
		#1		read = 32'd4022249759;
		#1		read = 32'd4032629328;
		#1		read = 32'd4042820384;
		#1		read = 32'd4052821908;
		#1		read = 32'd4062632899;
		#1		read = 32'd4072252378;
		#1		read = 32'd4081679381;
		#1		read = 32'd4090912966;
		#1		read = 32'd4099952210;
		#1		read = 32'd4108796208;
		#1		read = 32'd4117444077;
		#1		read = 32'd4125894951;
		#1		read = 32'd4134147986;
		#1		read = 32'd4142202357;
		#1		read = 32'd4150057257;
		#1		read = 32'd4157711901;
		#1		read = 32'd4165165524;
		#1		read = 32'd4172417381;
		#1		read = 32'd4179466746;
		#1		read = 32'd4186312914;
		#1		read = 32'd4192955201;
		#1		read = 32'd4199392943;
		#1		read = 32'd4205625495;
		#1		read = 32'd4211652235;
		#1		read = 32'd4217472560;
		#1		read = 32'd4223085888;
		#1		read = 32'd4228491657;
		#1		read = 32'd4233689327;
		#1		read = 32'd4238678379;
		#1		read = 32'd4243458312;
		#1		read = 32'd4248028650;
		#1		read = 32'd4252388935;
		#1		read = 32'd4256538732;
		#1		read = 32'd4260477624;
		#1		read = 32'd4264205219;
		#1		read = 32'd4267721144;
		#1		read = 32'd4271025046;
		#1		read = 32'd4274116596;
		#1		read = 32'd4276995485;
		#1		read = 32'd4279661424;
		#1		read = 32'd4282114148;
		#1		read = 32'd4284353410;
		#1		read = 32'd4286378986;
		#1		read = 32'd4288190675;
		#1		read = 32'd4289788296;
		#1		read = 32'd4291171687;
		#1		read = 32'd4292340711;
		#1		read = 32'd4293295252;
		#1		read = 32'd4294035213;
		#1		read = 32'd4294560521;
		#1		read = 32'd4294871123;
		#1		read = 32'd4294966988;
		#1		read = 32'd4294848106;
		#1		read = 32'd4294514490;
		#1		read = 32'd4293966172;
		#1		read = 32'd4293203208;
		#1		read = 32'd4292225674;
		#1		read = 32'd4291033667;
		#1		read = 32'd4289627307;
		#1		read = 32'd4288006735;
		#1		read = 32'd4286172112;
		#1		read = 32'd4284123622;
		#1		read = 32'd4281861470;
		#1		read = 32'd4279385882;
		#1		read = 32'd4276697105;
		#1		read = 32'd4273795409;
		#1		read = 32'd4270681083;
		#1		read = 32'd4267354439;
		#1		read = 32'd4263815810;
		#1		read = 32'd4260065550;
		#1		read = 32'd4256104033;
		#1		read = 32'd4251931656;
		#1		read = 32'd4247548836;
		#1		read = 32'd4242956011;
		#1		read = 32'd4238153641;
		#1		read = 32'd4233142205;
		#1		read = 32'd4227922205;
		#1		read = 32'd4222494163;
		#1		read = 32'd4216858622;
		#1		read = 32'd4211016145;
		#1		read = 32'd4204967316;
		#1		read = 32'd4198712741;
		#1		read = 32'd4192253045;
		#1		read = 32'd4185588873;
		#1		read = 32'd4178720893;
		#1		read = 32'd4171649790;
		#1		read = 32'd4164376273;
		#1		read = 32'd4156901068;
		#1		read = 32'd4149224923;
		#1		read = 32'd4141348605;
		#1		read = 32'd4133272903;
		#1		read = 32'd4124998623;
		#1		read = 32'd4116526594;
		#1		read = 32'd4107857662;
		#1		read = 32'd4098992694;
		#1		read = 32'd4089932577;
		#1		read = 32'd4080678216;
		#1		read = 32'd4071230538;
		#1		read = 32'd4061590487;
		#1		read = 32'd4051759026;
		#1		read = 32'd4041737140;
		#1		read = 32'd4031525830;
		#1		read = 32'd4021126117;
		#1		read = 32'd4010539041;
		#1		read = 32'd3999765662;
		#1		read = 32'd3988807056;
		#1		read = 32'd3977664319;
		#1		read = 32'd3966338565;
		#1		read = 32'd3954830928;
		#1		read = 32'd3943142557;
		#1		read = 32'd3931274622;
		#1		read = 32'd3919228309;
		#1		read = 32'd3907004823;
		#1		read = 32'd3894605387;
		#1		read = 32'd3882031240;
		#1		read = 32'd3869283640;
		#1		read = 32'd3856363861;
		#1		read = 32'd3843273195;
		#1		read = 32'd3830012952;
		#1		read = 32'd3816584457;
		#1		read = 32'd3802989054;
		#1		read = 32'd3789228102;
		#1		read = 32'd3775302976;
		#1		read = 32'd3761215070;
		#1		read = 32'd3746965792;
		#1		read = 32'd3732556567;
		#1		read = 32'd3717988836;
		#1		read = 32'd3703264056;
		#1		read = 32'd3688383700;
		#1		read = 32'd3673349254;
		#1		read = 32'd3658162224;
		#1		read = 32'd3642824126;
		#1		read = 32'd3627336496;
		#1		read = 32'd3611700882;
		#1		read = 32'd3595918847;
		#1		read = 32'd3579991970;
		#1		read = 32'd3563921844;
		#1		read = 32'd3547710074;
		#1		read = 32'd3531358283;
		#1		read = 32'd3514868106;
		#1		read = 32'd3498241192;
		#1		read = 32'd3481479203;
		#1		read = 32'd3464583816;
		#1		read = 32'd3447556719;
		#1		read = 32'd3430399617;
		#1		read = 32'd3413114223;
		#1		read = 32'd3395702268;
		#1		read = 32'd3378165492;
		#1		read = 32'd3360505649;
		#1		read = 32'd3342724505;
		#1		read = 32'd3324823838;
		#1		read = 32'd3306805437;
		#1		read = 32'd3288671106;
		#1		read = 32'd3270422656;
		#1		read = 32'd3252061914;
		#1		read = 32'd3233590714;
		#1		read = 32'd3215010905;
		#1		read = 32'd3196324344;
		#1		read = 32'd3177532900;
		#1		read = 32'd3158638452;
		#1		read = 32'd3139642889;
		#1		read = 32'd3120548111;
		#1		read = 32'd3101356028;
		#1		read = 32'd3082068558;
		#1		read = 32'd3062687630;
		#1		read = 32'd3043215183;
		#1		read = 32'd3023653163;
		#1		read = 32'd3004003527;
		#1		read = 32'd2984268240;
		#1		read = 32'd2964449275;
		#1		read = 32'd2944548614;
		#1		read = 32'd2924568247;
		#1		read = 32'd2904510172;
		#1		read = 32'd2884376396;
		#1		read = 32'd2864168931;
		#1		read = 32'd2843889797;
		#1		read = 32'd2823541024;
		#1		read = 32'd2803124646;
		#1		read = 32'd2782642704;
		#1		read = 32'd2762097247;
		#1		read = 32'd2741490329;
		#1		read = 32'd2720824010;
		#1		read = 32'd2700100358;
		#1		read = 32'd2679321445;
		#1		read = 32'd2658489349;
		#1		read = 32'd2637606152;
		#1		read = 32'd2616673944;
		#1		read = 32'd2595694817;
		#1		read = 32'd2574670869;
		#1		read = 32'd2553604203;
		#1		read = 32'd2532496925;
		#1		read = 32'd2511351146;
		#1		read = 32'd2490168981;
		#1		read = 32'd2468952547;
		#1		read = 32'd2447703967;
		#1		read = 32'd2426425365;
		#1		read = 32'd2405118869;
		#1		read = 32'd2383786610;
		#1		read = 32'd2362430720;
		#1		read = 32'd2341053337;
		#1		read = 32'd2319656596;
		#1		read = 32'd2298242638;
		#1		read = 32'd2276813605;
		#1		read = 32'd2255371638;
		#1		read = 32'd2233918883;
		#1		read = 32'd2212457484;
		#1		read = 32'd2190989588;
		#1		read = 32'd2169517342;
		#1		read = 32'd2148042892;
		#1		read = 32'd2126568386;
		#1		read = 32'd2105095972;
		#1		read = 32'd2083627796;
		#1		read = 32'd2062166006;
		#1		read = 32'd2040712748;
		#1		read = 32'd2019270166;
		#1		read = 32'd1997840406;
		#1		read = 32'd1976425610;
		#1		read = 32'd1955027920;
		#1		read = 32'd1933649475;
		#1		read = 32'd1912292414;
		#1		read = 32'd1890958871;
		#1		read = 32'd1869650981;
		#1		read = 32'd1848370873;
		#1		read = 32'd1827120677;
		#1		read = 32'd1805902517;
		#1		read = 32'd1784718514;
		#1		read = 32'd1763570788;
		#1		read = 32'd1742461453;
		#1		read = 32'd1721392619;
		#1		read = 32'd1700366395;
		#1		read = 32'd1679384881;
		#1		read = 32'd1658450178;
		#1		read = 32'd1637564377;
		#1		read = 32'd1616729567;
		#1		read = 32'd1595947833;
		#1		read = 32'd1575221252;
		#1		read = 32'd1554551896;
		#1		read = 32'd1533941833;
		#1		read = 32'd1513393124;
		#1		read = 32'd1492907823;
		#1		read = 32'd1472487980;
		#1		read = 32'd1452135635;
		#1		read = 32'd1431852825;
		#1		read = 32'd1411641577;
		#1		read = 32'd1391503913;
		#1		read = 32'd1371441846;
		#1		read = 32'd1351457382;
		#1		read = 32'd1331552521;
		#1		read = 32'd1311729252;
		#1		read = 32'd1291989557;
		#1		read = 32'd1272335412;
		#1		read = 32'd1252768780;
		#1		read = 32'd1233291620;
		#1		read = 32'd1213905877;
		#1		read = 32'd1194613492;
		#1		read = 32'd1175416393;
		#1		read = 32'd1156316500;
		#1		read = 32'd1137315722;
		#1		read = 32'd1118415961;
		#1		read = 32'd1099619106;
		#1		read = 32'd1080927036;
		#1		read = 32'd1062341621;
		#1		read = 32'd1043864719;
		#1		read = 32'd1025498178;
		#1		read = 32'd1007243835;
		#1		read = 32'd989103515;
		#1		read = 32'd971079032;
		#1		read = 32'd953172188;
		#1		read = 32'd935384774;
		#1		read = 32'd917718570;
		#1		read = 32'd900175341;
		#1		read = 32'd882756841;
		#1		read = 32'd865464814;
		#1		read = 32'd848300987;
		#1		read = 32'd831267077;
		#1		read = 32'd814364788;
		#1		read = 32'd797595809;
		#1		read = 32'd780961819;
		#1		read = 32'd764464479;
		#1		read = 32'd748105440;
		#1		read = 32'd731886338;
		#1		read = 32'd715808794;
		#1		read = 32'd699874417;
		#1		read = 32'd684084799;
		#1		read = 32'd668441520;
		#1		read = 32'd652946144;
		#1		read = 32'd637600221;
		#1		read = 32'd622405284;
		#1		read = 32'd607362854;
		#1		read = 32'd592474435;
		#1		read = 32'd577741516;
		#1		read = 32'd563165569;
		#1		read = 32'd548748053;
		#1		read = 32'd534490409;
		#1		read = 32'd520394063;
		#1		read = 32'd506460425;
		#1		read = 32'd492690888;
		#1		read = 32'd479086828;
		#1		read = 32'd465649607;
		#1		read = 32'd452380568;
		#1		read = 32'd439281038;
		#1		read = 32'd426352326;
		#1		read = 32'd413595727;
		#1		read = 32'd401012514;
		#1		read = 32'd388603948;
		#1		read = 32'd376371267;
		#1		read = 32'd364315697;
		#1		read = 32'd352438442;
		#1		read = 32'd340740690;
		#1		read = 32'd329223611;
		#1		read = 32'd317888356;
		#1		read = 32'd306736059;
		#1		read = 32'd295767835;
		#1		read = 32'd284984782;
		#1		read = 32'd274387977;
		#1		read = 32'd263978479;
		#1		read = 32'd253757331;
		#1		read = 32'd243725554;
		#1		read = 32'd233884151;
		#1		read = 32'd224234106;
		#1		read = 32'd214776385;
		#1		read = 32'd205511933;
		#1		read = 32'd196441676;
		#1		read = 32'd187566522;
		#1		read = 32'd178887358;
		#1		read = 32'd170405052;
		#1		read = 32'd162120453;
		#1		read = 32'd154034388;
		#1		read = 32'd146147666;
		#1		read = 32'd138461076;
		#1		read = 32'd130975387;
		#1		read = 32'd123691346;
		#1		read = 32'd116609684;
		#1		read = 32'd109731107;
		#1		read = 32'd103056304;
		#1		read = 32'd96585941;
		#1		read = 32'd90320667;
		#1		read = 32'd84261107;
		#1		read = 32'd78407868;
		#1		read = 32'd72761535;
		#1		read = 32'd67322672;
		#1		read = 32'd62091824;
		#1		read = 32'd57069513;
		#1		read = 32'd52256241;
		#1		read = 32'd47652491;
		#1		read = 32'd43258722;
		#1		read = 32'd39075374;
		#1		read = 32'd35102865;
		#1		read = 32'd31341592;
		#1		read = 32'd27791931;
		#1		read = 32'd24454238;
		#1		read = 32'd21328847;
		#1		read = 32'd18416068;
		#1		read = 32'd15716195;
		#1		read = 32'd13229497;
		#1		read = 32'd10956223;
		#1		read = 32'd8896599;
		#1		read = 32'd7050832;
		#1		read = 32'd5419107;
		#1		read = 32'd4001587;
		#1		read = 32'd2798413;
		#1		read = 32'd1809705;
		#1		read = 32'd1035564;
		#1		read = 32'd476065;
		#1		read = 32'd131265;
		#1		read = 32'd1199;
		#1		read = 32'd85879;
		#1		read = 32'd385297;
		#1		read = 32'd899424;
		#1		read = 32'd1628206;
		#1		read = 32'd2571573;
		#1		read = 32'd3729429;
		#1		read = 32'd5101659;
		#1		read = 32'd6688125;
		#1		read = 32'd8488669;
		#1		read = 32'd10503110;
		#1		read = 32'd12731248;
		#1		read = 32'd15172859;
		#1		read = 32'd17827700;
		#1		read = 32'd20695504;
		#1		read = 32'd23775986;
		#1		read = 32'd27068836;
		#1		read = 32'd30573726;
		#1		read = 32'd34290306;
		#1		read = 32'd38218203;
		#1		read = 32'd42357025;
		#1		read = 32'd46706357;
		#1		read = 32'd51265766;
		#1		read = 32'd56034795;
		#1		read = 32'd61012966;
		#1		read = 32'd66199784;
		#1		read = 32'd71594727;
		#1		read = 32'd77197258;
		#1		read = 32'd83006816;
		#1		read = 32'd89022820;
		#1		read = 32'd95244668;
		#1		read = 32'd101671739;
		#1		read = 32'd108303389;
		#1		read = 32'd115138955;
		#1		read = 32'd122177754;
		#1		read = 32'd129419082;
		#1		read = 32'd136862214;
		#1		read = 32'd144506407;
		#1		read = 32'd152350897;
		#1		read = 32'd160394897;
		#1		read = 32'd168637606;
		#1		read = 32'd177078196;
		#1		read = 32'd185715826;
		#1		read = 32'd194549631;
		#1		read = 32'd203578728;
		#1		read = 32'd212802214;
		#1		read = 32'd222219166;
		#1		read = 32'd231828643;
		#1		read = 32'd241629684;
		#1		read = 32'd251621309;
		#1		read = 32'd261802518;
		#1		read = 32'd272172294;
		#1		read = 32'd282729600;
		#1		read = 32'd293473379;
		#1		read = 32'd304402558;
		#1		read = 32'd315516043;
		#1		read = 32'd326812724;
		#1		read = 32'd338291470;
		#1		read = 32'd349951134;
		#1		read = 32'd361790550;
		#1		read = 32'd373808534;
		#1		read = 32'd386003883;
		#1		read = 32'd398375379;
		#1		read = 32'd410921785;
		#1		read = 32'd423641845;
		#1		read = 32'd436534288;
		#1		read = 32'd449597824;
		#1		read = 32'd462831148;
		#1		read = 32'd476232935;
		#1		read = 32'd489801846;
		#1		read = 32'd503536524;
		#1		read = 32'd517435595;
		#1		read = 32'd531497670;
		#1		read = 32'd545721342;
		#1		read = 32'd560105189;
		#1		read = 32'd574647772;
		#1		read = 32'd589347638;
		#1		read = 32'd604203316;
		#1		read = 32'd619213321;
		#1		read = 32'd634376151;
		#1		read = 32'd649690291;
		#1		read = 32'd665154209;
		#1		read = 32'd680766359;
		#1		read = 32'd696525179;
		#1		read = 32'd712429094;
		#1		read = 32'd728476513;
		#1		read = 32'd744665832;
		#1		read = 32'd760995431;
		#1		read = 32'd777463678;
		#1		read = 32'd794068926;
		#1		read = 32'd810809514;
		#1		read = 32'd827683769;
		#1		read = 32'd844690002;
		#1		read = 32'd861826514;
		#1		read = 32'd879091590;
		#1		read = 32'd896483504;
		#1		read = 32'd914000518;
		#1		read = 32'd931640878;
		#1		read = 32'd949402822;
		#1		read = 32'd967284573;
		#1		read = 32'd985284343;
		#1		read = 32'd1003400332;
		#1		read = 32'd1021630729;
		#1		read = 32'd1039973709;
		#1		read = 32'd1058427440;
		#1		read = 32'd1076990075;
		#1		read = 32'd1095659759;
		#1		read = 32'd1114434625;
		#1		read = 32'd1133312794;
		#1		read = 32'd1152292380;
		#1		read = 32'd1171371484;
		#1		read = 32'd1190548198;
		#1		read = 32'd1209820605;
		#1		read = 32'd1229186778;
		#1		read = 32'd1248644780;
		#1		read = 32'd1268192664;
		#1		read = 32'd1287828477;
		#1		read = 32'd1307550255;
		#1		read = 32'd1327356026;
		#1		read = 32'd1347243808;
		#1		read = 32'd1367211614;
		#1		read = 32'd1387257447;
		#1		read = 32'd1407379301;
		#1		read = 32'd1427575166;
		#1		read = 32'd1447843020;
		#1		read = 32'd1468180838;
		#1		read = 32'd1488586586;
		#1		read = 32'd1509058223;
		#1		read = 32'd1529593702;
		#1		read = 32'd1550190969;
		#1		read = 32'd1570847965;
		#1		read = 32'd1591562624;
		#1		read = 32'd1612332875;
		#1		read = 32'd1633156641;
		#1		read = 32'd1654031839;
		#1		read = 32'd1674956381;
		#1		read = 32'd1695928176;
		#1		read = 32'd1716945126;
		#1		read = 32'd1738005130;
		#1		read = 32'd1759106081;
		#1		read = 32'd1780245869;
		#1		read = 32'd1801422381;
		#1		read = 32'd1822633499;
		#1		read = 32'd1843877101;
		#1		read = 32'd1865151064;
		#1		read = 32'd1886453260;
		#1		read = 32'd1907781559;
		#1		read = 32'd1929133828;
		#1		read = 32'd1950507931;
		#1		read = 32'd1971901732;
		#1		read = 32'd1993313091;
		#1		read = 32'd2014739867;
		#1		read = 32'd2036179918;
		#1		read = 32'd2057631098;
		#1		read = 32'd2079091264;
		#1		read = 32'd2100558269;
		#1		read = 32'd2122029966;
		#1		read = 32'd2143504209;
		#1		read = 32'd2164978850;
		#1		read = 32'd2186451741;
		#1		read = 32'd2207920735;
		#1		read = 32'd2229383686;
		#1		read = 32'd2250838447;
		#1		read = 32'd2272282872;
		#1		read = 32'd2293714818;
		#1		read = 32'd2315132140;
		#1		read = 32'd2336532698;
		#1		read = 32'd2357914351;
		#1		read = 32'd2379274961;
		#1		read = 32'd2400612393;
		#1		read = 32'd2421924511;
		#1		read = 32'd2443209186;
		#1		read = 32'd2464464289;
		#1		read = 32'd2485687693;
		#1		read = 32'd2506877278;
		#1		read = 32'd2528030923;
		#1		read = 32'd2549146514;
		#1		read = 32'd2570221939;
		#1		read = 32'd2591255091;
		#1		read = 32'd2612243866;
		#1		read = 32'd2633186165;
		#1		read = 32'd2654079895;
		#1		read = 32'd2674922965;
		#1		read = 32'd2695713291;
		#1		read = 32'd2716448796;
		#1		read = 32'd2737127404;
		#1		read = 32'd2757747048;
		#1		read = 32'd2778305666;
		#1		read = 32'd2798801203;
		#1		read = 32'd2819231609;
		#1		read = 32'd2839594840;
		#1		read = 32'd2859888861;
		#1		read = 32'd2880111642;
		#1		read = 32'd2900261160;
		#1		read = 32'd2920335402;
		#1		read = 32'd2940332359;
		#1		read = 32'd2960250032;
		#1		read = 32'd2980086428;
		#1		read = 32'd2999839566;
		#1		read = 32'd3019507468;
		#1		read = 32'd3039088169;
		#1		read = 32'd3058579710;
		#1		read = 32'd3077980142;
		#1		read = 32'd3097287525;
		#1		read = 32'd3116499929;
		#1		read = 32'd3135615432;
		#1		read = 32'd3154632122;
		#1		read = 32'd3173548099;
		#1		read = 32'd3192361469;
		#1		read = 32'd3211070353;
		#1		read = 32'd3229672880;
		#1		read = 32'd3248167188;
		#1		read = 32'd3266551429;
		#1		read = 32'd3284823763;
		#1		read = 32'd3302982365;
		#1		read = 32'd3321025418;
		#1		read = 32'd3338951118;
		#1		read = 32'd3356757672;
		#1		read = 32'd3374443299;
		#1		read = 32'd3392006232;
		#1		read = 32'd3409444713;
		#1		read = 32'd3426757000;
		#1		read = 32'd3443941360;
		#1		read = 32'd3460996075;
		#1		read = 32'd3477919441;
		#1		read = 32'd3494709763;
		#1		read = 32'd3511365365;
		#1		read = 32'd3527884579;
		#1		read = 32'd3544265754;
		#1		read = 32'd3560507252;
		#1		read = 32'd3576607450;
		#1		read = 32'd3592564735;
		#1		read = 32'd3608377514;
		#1		read = 32'd3624044205;
		#1		read = 32'd3639563241;
		#1		read = 32'd3654933071;
		#1		read = 32'd3670152156;
		#1		read = 32'd3685218976;
		#1		read = 32'd3700132024;
		#1		read = 32'd3714889808;
		#1		read = 32'd3729490853;
		#1		read = 32'd3743933698;
		#1		read = 32'd3758216900;
		#1		read = 32'd3772339030;
		#1		read = 32'd3786298676;
		#1		read = 32'd3800094441;
		#1		read = 32'd3813724947;
		#1		read = 32'd3827188830;
		#1		read = 32'd3840484744;
		#1		read = 32'd3853611359;
		#1		read = 32'd3866567363;
		#1		read = 32'd3879351460;
		#1		read = 32'd3891962372;
		#1		read = 32'd3904398837;
		#1		read = 32'd3916659612;
		#1		read = 32'd3928743471;
		#1		read = 32'd3940649206;
		#1		read = 32'd3952375625;
		#1		read = 32'd3963921557;
		#1		read = 32'd3975285847;
		#1		read = 32'd3986467358;
		#1		read = 32'd3997464972;
		#1		read = 32'd4008277589;
		#1		read = 32'd4018904128;
		#1		read = 32'd4029343527;
		#1		read = 32'd4039594742;
		#1		read = 32'd4049656747;
		#1		read = 32'd4059528537;
		#1		read = 32'd4069209123;
		#1		read = 32'd4078697539;
		#1		read = 32'd4087992834;
		#1		read = 32'd4097094081;
		#1		read = 32'd4106000368;
		#1		read = 32'd4114710805;
		#1		read = 32'd4123224521;
		#1		read = 32'd4131540664;
		#1		read = 32'd4139658404;
		#1		read = 32'd4147576927;
		#1		read = 32'd4155295443;
		#1		read = 32'd4162813180;
		#1		read = 32'd4170129385;
		#1		read = 32'd4177243327;
		#1		read = 32'd4184154295;
		#1		read = 32'd4190861598;
		#1		read = 32'd4197364564;
		#1		read = 32'd4203662544;
		#1		read = 32'd4209754908;
		#1		read = 32'd4215641047;
		#1		read = 32'd4221320372;
		#1		read = 32'd4226792314;
		#1		read = 32'd4232056328;
		#1		read = 32'd4237111886;
		#1		read = 32'd4241958483;
		#1		read = 32'd4246595634;
		#1		read = 32'd4251022875;
		#1		read = 32'd4255239765;
		#1		read = 32'd4259245881;
		#1		read = 32'd4263040822;
		#1		read = 32'd4266624209;
		#1		read = 32'd4269995684;
		#1		read = 32'd4273154909;
		#1		read = 32'd4276101570;
		#1		read = 32'd4278835370;
		#1		read = 32'd4281356036;
		#1		read = 32'd4283663318;
		#1		read = 32'd4285756983;
		#1		read = 32'd4287636822;
		#1		read = 32'd4289302648;
		#1		read = 32'd4290754294;
		#1		read = 32'd4291991615;
		#1		read = 32'd4293014487;
		#1		read = 32'd4293822807;
		#1		read = 32'd4294416495;
		#1		read = 32'd4294795492;
		#1		read = 32'd4294959759;
		#1		read = 32'd4294909281;
		#1		read = 32'd4294644061;
		#1		read = 32'd4294164128;
		#1		read = 32'd4293469528;
		#1		read = 32'd4292560331;
		#1		read = 32'd4291436629;
		#1		read = 32'd4290098533;
		#1		read = 32'd4288546177;
		#1		read = 32'd4286779717;
		#1		read = 32'd4284799329;
		#1		read = 32'd4282605211;
		#1		read = 32'd4280197583;
		#1		read = 32'd4277576685;
		#1		read = 32'd4274742780;
		#1		read = 32'd4271696150;
		#1		read = 32'd4268437102;
		#1		read = 32'd4264965959;
		#1		read = 32'd4261283070;
		#1		read = 32'd4257388803;
		#1		read = 32'd4253283547;
		#1		read = 32'd4248967713;
		#1		read = 32'd4244441732;
		#1		read = 32'd4239706057;
		#1		read = 32'd4234761162;
		#1		read = 32'd4229607540;
		#1		read = 32'd4224245708;
		#1		read = 32'd4218676202;
		#1		read = 32'd4212899578;
		#1		read = 32'd4206916414;
		#1		read = 32'd4200727309;
		#1		read = 32'd4194332880;
		#1		read = 32'd4187733769;
		#1		read = 32'd4180930634;
		#1		read = 32'd4173924157;
		#1		read = 32'd4166715037;
		#1		read = 32'd4159303995;
		#1		read = 32'd4151691774;
		#1		read = 32'd4143879133;
		#1		read = 32'd4135866854;
		#1		read = 32'd4127655738;
		#1		read = 32'd4119246607;
		#1		read = 32'd4110640301;
		#1		read = 32'd4101837682;
		#1		read = 32'd4092839628;
		#1		read = 32'd4083647041;
		#1		read = 32'd4074260838;
		#1		read = 32'd4064681960;
		#1		read = 32'd4054911363;
		#1		read = 32'd4044950026;
		#1		read = 32'd4034798943;
		#1		read = 32'd4024459130;
		#1		read = 32'd4013931621;
		#1		read = 32'd4003217469;
		#1		read = 32'd3992317745;
		#1		read = 32'd3981233540;
		#1		read = 32'd3969965961;
		#1		read = 32'd3958516135;
		#1		read = 32'd3946885207;
		#1		read = 32'd3935074341;
		#1		read = 32'd3923084717;
		#1		read = 32'd3910917534;
		#1		read = 32'd3898574010;
		#1		read = 32'd3886055378;
		#1		read = 32'd3873362890;
		#1		read = 32'd3860497816;
		#1		read = 32'd3847461442;
		#1		read = 32'd3834255071;
		#1		read = 32'd3820880025;
		#1		read = 32'd3807337641;
		#1		read = 32'd3793629272;
		#1		read = 32'd3779756290;
		#1		read = 32'd3765720083;
		#1		read = 32'd3751522053;
		#1		read = 32'd3737163620;
		#1		read = 32'd3722646221;
		#1		read = 32'd3707971307;
		#1		read = 32'd3693140346;
		#1		read = 32'd3678154820;
		#1		read = 32'd3663016228;
		#1		read = 32'd3647726084;
		#1		read = 32'd3632285918;
		#1		read = 32'd3616697272;
		#1		read = 32'd3600961706;
		#1		read = 32'd3585080793;
		#1		read = 32'd3569056123;
		#1		read = 32'd3552889295;
		#1		read = 32'd3536581929;
		#1		read = 32'd3520135654;
		#1		read = 32'd3503552115;
		#1		read = 32'd3486832970;
		#1		read = 32'd3469979891;
		#1		read = 32'd3452994564;
		#1		read = 32'd3435878687;
		#1		read = 32'd3418633971;
		#1		read = 32'd3401262142;
		#1		read = 32'd3383764935;
		#1		read = 32'd3366144102;
		#1		read = 32'd3348401403;
		#1		read = 32'd3330538614;
		#1		read = 32'd3312557520;
		#1		read = 32'd3294459920;
		#1		read = 32'd3276247623;
		#1		read = 32'd3257922450;
		#1		read = 32'd3239486235;
		#1		read = 32'd3220940820;
		#1		read = 32'd3202288061;
		#1		read = 32'd3183529822;
		#1		read = 32'd3164667979;
		#1		read = 32'd3145704419;
		#1		read = 32'd3126641037;
		#1		read = 32'd3107479740;
		#1		read = 32'd3088222445;
		#1		read = 32'd3068871077;
		#1		read = 32'd3049427570;
		#1		read = 32'd3029893870;
		#1		read = 32'd3010271930;
		#1		read = 32'd2990563711;
		#1		read = 32'd2970771185;
		#1		read = 32'd2950896331;
		#1		read = 32'd2930941137;
		#1		read = 32'd2910907597;
		#1		read = 32'd2890797716;
		#1		read = 32'd2870613504;
		#1		read = 32'd2850356980;
		#1		read = 32'd2830030168;
		#1		read = 32'd2809635103;
		#1		read = 32'd2789173823;
		#1		read = 32'd2768648375;
		#1		read = 32'd2748060810;
		#1		read = 32'd2727413189;
		#1		read = 32'd2706707575;
		#1		read = 32'd2685946039;
		#1		read = 32'd2665130657;
		#1		read = 32'd2644263511;
		#1		read = 32'd2623346687;
		#1		read = 32'd2602382278;
		#1		read = 32'd2581372379;
		#1		read = 32'd2560319091;
		#1		read = 32'd2539224521;
		#1		read = 32'd2518090776;
		#1		read = 32'd2496919971;
		#1		read = 32'd2475714223;
		#1		read = 32'd2454475652;
		#1		read = 32'd2433206382;
		#1		read = 32'd2411908540;
		#1		read = 32'd2390584256;
		#1		read = 32'd2369235662;
		#1		read = 32'd2347864893;
		#1		read = 32'd2326474086;
		#1		read = 32'd2305065380;
		#1		read = 32'd2283640916;
		#1		read = 32'd2262202836;
		#1		read = 32'd2240753285;
		#1		read = 32'd2219294406;
		#1		read = 32'd2197828347;
		#1		read = 32'd2176357253;
		#1		read = 32'd2154883272;
		#1		read = 32'd2133408551;
		#1		read = 32'd2111935238;
		#1		read = 32'd2090465479;
		#1		read = 32'd2069001422;
		#1		read = 32'd2047545213;
		#1		read = 32'd2026098998;
		#1		read = 32'd2004664921;
		#1		read = 32'd1983245126;
		#1		read = 32'd1961841755;
		#1		read = 32'd1940456948;
		#1		read = 32'd1919092843;
		#1		read = 32'd1897751577;
		#1		read = 32'd1876435285;
		#1		read = 32'd1855146096;
		#1		read = 32'd1833886142;
		#1		read = 32'd1812657547;
		#1		read = 32'd1791462434;
		#1		read = 32'd1770302923;
		#1		read = 32'd1749181129;
		#1		read = 32'd1728099166;
		#1		read = 32'd1707059141;
		#1		read = 32'd1686063157;
		#1		read = 32'd1665113316;
		#1		read = 32'd1644211711;
		#1		read = 32'd1623360433;
		#1		read = 32'd1602561567;
		#1		read = 32'd1581817192;
		#1		read = 32'd1561129384;
		#1		read = 32'd1540500211;
		#1		read = 32'd1519931735;
		#1		read = 32'd1499426014;
		#1		read = 32'd1478985099;
		#1		read = 32'd1458611032;
		#1		read = 32'd1438305853;
		#1		read = 32'd1418071590;
		#1		read = 32'd1397910268;
		#1		read = 32'd1377823903;
		#1		read = 32'd1357814503;
		#1		read = 32'd1337884070;
		#1		read = 32'd1318034595;
		#1		read = 32'd1298268065;
		#1		read = 32'd1278586456;
		#1		read = 32'd1258991736;
		#1		read = 32'd1239485864;
		#1		read = 32'd1220070791;
		#1		read = 32'd1200748459;
		#1		read = 32'd1181520800;
		#1		read = 32'd1162389736;
		#1		read = 32'd1143357180;
		#1		read = 32'd1124425037;
		#1		read = 32'd1105595198;
		#1		read = 32'd1086869547;
		#1		read = 32'd1068249957;
		#1		read = 32'd1049738290;
		#1		read = 32'd1031336396;
		#1		read = 32'd1013046115;
		#1		read = 32'd994869278;
		#1		read = 32'd976807701;
		#1		read = 32'd958863191;
		#1		read = 32'd941037541;
		#1		read = 32'd923332536;
		#1		read = 32'd905749944;
		#1		read = 32'd888291525;
		#1		read = 32'd870959024;
		#1		read = 32'd853754174;
		#1		read = 32'd836678696;
		#1		read = 32'd819734298;
		#1		read = 32'd802922673;
		#1		read = 32'd786245503;
		#1		read = 32'd769704457;
		#1		read = 32'd753301186;
		#1		read = 32'd737037333;
		#1		read = 32'd720914524;
		#1		read = 32'd704934370;
		#1		read = 32'd689098470;
		#1		read = 32'd673408407;
		#1		read = 32'd657865750;
		#1		read = 32'd642472054;
		#1		read = 32'd627228858;
		#1		read = 32'd612137686;
		#1		read = 32'd597200048;
		#1		read = 32'd582417436;
		#1		read = 32'd567791330;
		#1		read = 32'd553323192;
		#1		read = 32'd539014468;
		#1		read = 32'd524866590;
		#1		read = 32'd510880972;
		#1		read = 32'd497059014;
		#1		read = 32'd483402096;
		#1		read = 32'd469911585;
		#1		read = 32'd456588830;
		#1		read = 32'd443435163;
		#1		read = 32'd430451899;
		#1		read = 32'd417640338;
		#1		read = 32'd405001759;
		#1		read = 32'd392537426;
		#1		read = 32'd380248587;
		#1		read = 32'd368136470;
		#1		read = 32'd356202287;
		#1		read = 32'd344447229;
		#1		read = 32'd332872474;
		#1		read = 32'd321479179;
		#1		read = 32'd310268483;
		#1		read = 32'd299241506;
		#1		read = 32'd288399352;
		#1		read = 32'd277743105;
		#1		read = 32'd267273831;
		#1		read = 32'd256992576;
		#1		read = 32'd246900368;
		#1		read = 32'd236998218;
		#1		read = 32'd227287114;
		#1		read = 32'd217768028;
		#1		read = 32'd208441912;
		#1		read = 32'd199309699;
		#1		read = 32'd190372302;
		#1		read = 32'd181630614;
		#1		read = 32'd173085510;
		#1		read = 32'd164737843;
		#1		read = 32'd156588450;
		#1		read = 32'd148638145;
		#1		read = 32'd140887723;
		#1		read = 32'd133337958;
		#1		read = 32'd125989606;
		#1		read = 32'd118843402;
		#1		read = 32'd111900061;
		#1		read = 32'd105160276;
		#1		read = 32'd98624722;
		#1		read = 32'd92294052;
		#1		read = 32'd86168899;
		#1		read = 32'd80249876;
		#1		read = 32'd74537574;
		#1		read = 32'd69032566;
		#1		read = 32'd63735401;
		#1		read = 32'd58646608;
		#1		read = 32'd53766698;
		#1		read = 32'd49096158;
		#1		read = 32'd44635455;
		#1		read = 32'd40385035;
		#1		read = 32'd36345323;
		#1		read = 32'd32516723;
		#1		read = 32'd28899618;
		#1		read = 32'd25494370;
		#1		read = 32'd22301318;
		#1		read = 32'd19320784;
		#1		read = 32'd16553063;
		#1		read = 32'd13998435;
		#1		read = 32'd11657152;
		#1		read = 32'd9529451;
		#1		read = 32'd7615543;
		#1		read = 32'd5915621;
		#1		read = 32'd4429853;
		#1		read = 32'd3158389;
		#1		read = 32'd2101356;
		#1		read = 32'd1258859;
		#1		read = 32'd630983;
		#1		read = 32'd217790;
		#1		read = 32'd19322;
		#1		read = 32'd35599;
		#1		read = 32'd266618;
		#1		read = 32'd712358;
		#1		read = 32'd1372773;
		#1		read = 32'd2247797;
		#1		read = 32'd3337344;
		#1		read = 32'd4641302;
		#1		read = 32'd6159544;
		#1		read = 32'd7891916;
		#1		read = 32'd9838245;
		#1		read = 32'd11998337;
		#1		read = 32'd14371976;
		#1		read = 32'd16958925;
		#1		read = 32'd19758924;
		#1		read = 32'd22771693;
		#1		read = 32'd25996933;
		#1		read = 32'd29434319;
		#1		read = 32'd33083508;
		#1		read = 32'd36944135;
		#1		read = 32'd41015815;
		#1		read = 32'd45298140;
		#1		read = 32'd49790681;
		#1		read = 32'd54492990;
		#1		read = 32'd59404596;
		#1		read = 32'd64525009;
		#1		read = 32'd69853716;
		#1		read = 32'd75390183;
		#1		read = 32'd81133859;
		#1		read = 32'd87084168;
		#1		read = 32'd93240515;
		#1		read = 32'd99602284;
		#1		read = 32'd106168840;
		#1		read = 32'd112939526;
		#1		read = 32'd119913665;
		#1		read = 32'd127090559;
		#1		read = 32'd134469490;
		#1		read = 32'd142049721;
		#1		read = 32'd149830494;
		#1		read = 32'd157811031;
		#1		read = 32'd165990533;
		#1		read = 32'd174368183;
		#1		read = 32'd182943143;
		#1		read = 32'd191714555;
		#1		read = 32'd200681542;
		#1		read = 32'd209843208;
		#1		read = 32'd219198637;
		#1		read = 32'd228746892;
		#1		read = 32'd238487019;
		#1		read = 32'd248418045;
		#1		read = 32'd258538975;
		#1		read = 32'd268848799;
		#1		read = 32'd279346484;
		#1		read = 32'd290030981;
		#1		read = 32'd300901223;
		#1		read = 32'd311956121;
		#1		read = 32'd323194570;
		#1		read = 32'd334615446;
		#1		read = 32'd346217608;
		#1		read = 32'd357999895;
		#1		read = 32'd369961129;
		#1		read = 32'd382100113;
		#1		read = 32'd394415635;
		#1		read = 32'd406906461;
		#1		read = 32'd419571344;
		#1		read = 32'd432409017;
		#1		read = 32'd445418196;
		#1		read = 32'd458597580;
		#1		read = 32'd471945851;
		#1		read = 32'd485461675;
		#1		read = 32'd499143699;
		#1		read = 32'd512990556;
		#1		read = 32'd527000861;
		#1		read = 32'd541173213;
		#1		read = 32'd555506195;
		#1		read = 32'd569998373;
		#1		read = 32'd584648298;
		#1		read = 32'd599454505;
		#1		read = 32'd614415514;
		#1		read = 32'd629529829;
		#1		read = 32'd644795938;
		#1		read = 32'd660212314;
		#1		read = 32'd675777416;
		#1		read = 32'd691489688;
		#1		read = 32'd707347557;
		#1		read = 32'd723349440;
		#1		read = 32'd739493734;
		#1		read = 32'd755778826;
		#1		read = 32'd772203088;
		#1		read = 32'd788764876;
		#1		read = 32'd805462535;
		#1		read = 32'd822294395;
		#1		read = 32'd839258773;
		#1		read = 32'd856353973;
		#1		read = 32'd873578284;
		#1		read = 32'd890929985;
		#1		read = 32'd908407340;
		#1		read = 32'd926008601;
		#1		read = 32'd943732010;
		#1		read = 32'd961575792;
		#1		read = 32'd979538164;
		#1		read = 32'd997617330;
		#1		read = 32'd1015811481;
		#1		read = 32'd1034118799;
		#1		read = 32'd1052537452;
		#1		read = 32'd1071065599;
		#1		read = 32'd1089701386;
		#1		read = 32'd1108442952;
		#1		read = 32'd1127288420;
		#1		read = 32'd1146235907;
		#1		read = 32'd1165283518;
		#1		read = 32'd1184429348;
		#1		read = 32'd1203671483;
		#1		read = 32'd1223007998;
		#1		read = 32'd1242436960;
		#1		read = 32'd1261956426;
		#1		read = 32'd1281564444;
		#1		read = 32'd1301259053;
		#1		read = 32'd1321038284;
		#1		read = 32'd1340900158;
		#1		read = 32'd1360842691;
		#1		read = 32'd1380863887;
		#1		read = 32'd1400961744;
		#1		read = 32'd1421134253;
		#1		read = 32'd1441379396;
		#1		read = 32'd1461695149;
		#1		read = 32'd1482079480;
		#1		read = 32'd1502530351;
		#1		read = 32'd1523045717;
		#1		read = 32'd1543623526;
		#1		read = 32'd1564261720;
		#1		read = 32'd1584958237;
		#1		read = 32'd1605711005;
		#1		read = 32'd1626517950;
		#1		read = 32'd1647376992;
		#1		read = 32'd1668286043;
		#1		read = 32'd1689243014;
		#1		read = 32'd1710245809;
		#1		read = 32'd1731292327;
		#1		read = 32'd1752380464;
		#1		read = 32'd1773508110;
		#1		read = 32'd1794673154;
		#1		read = 32'd1815873479;
		#1		read = 32'd1837106965;
		#1		read = 32'd1858371488;
		#1		read = 32'd1879664922;
		#1		read = 32'd1900985137;
		#1		read = 32'd1922330003;
		#1		read = 32'd1943697383;
		#1		read = 32'd1965085142;
		#1		read = 32'd1986491140;
		#1		read = 32'd2007913238;
		#1		read = 32'd2029349293;
		#1		read = 32'd2050797161;
		#1		read = 32'd2072254697;
		#1		read = 32'd2093719757;
		#1		read = 32'd2115190192;
		#1		read = 32'd2136663857;
		#1		read = 32'd2158138604;
		#1		read = 32'd2179612286;
		#1		read = 32'd2201082754;
		#1		read = 32'd2222547863;
		#1		read = 32'd2244005466;
		#1		read = 32'd2265453416;
		#1		read = 32'd2286889569;
		#1		read = 32'd2308311782;
		#1		read = 32'd2329717913;
		#1		read = 32'd2351105820;
		#1		read = 32'd2372473365;
		#1		read = 32'd2393818411;
		#1		read = 32'd2415138824;
		#1		read = 32'd2436432472;
		#1		read = 32'd2457697225;
		#1		read = 32'd2478930956;
		#1		read = 32'd2500131544;
		#1		read = 32'd2521296867;
		#1		read = 32'd2542424809;
		#1		read = 32'd2563513257;
		#1		read = 32'd2584560102;
		#1		read = 32'd2605563241;
		#1		read = 32'd2626520571;
		#1		read = 32'd2647429999;
		#1		read = 32'd2668289432;
		#1		read = 32'd2689096785;
		#1		read = 32'd2709849977;
		#1		read = 32'd2730546933;
		#1		read = 32'd2751185583;
		#1		read = 32'd2771763864;
		#1		read = 32'd2792279717;
		#1		read = 32'd2812731090;
		#1		read = 32'd2833115940;
		#1		read = 32'd2853432227;
		#1		read = 32'd2873677920;
		#1		read = 32'd2893850994;
		#1		read = 32'd2913949432;
		#1		read = 32'd2933971224;
		#1		read = 32'd2953914367;
		#1		read = 32'd2973776869;
		#1		read = 32'd2993556741;
		#1		read = 32'd3013252008;
		#1		read = 32'd3032860698;
		#1		read = 32'd3052380851;
		#1		read = 32'd3071810515;
		#1		read = 32'd3091147747;
		#1		read = 32'd3110390614;
		#1		read = 32'd3129537190;
		#1		read = 32'd3148585562;
		#1		read = 32'd3167533825;
		#1		read = 32'd3186380084;
		#1		read = 32'd3205122454;
		#1		read = 32'd3223759060;
		#1		read = 32'd3242288041;
		#1		read = 32'd3260707541;
		#1		read = 32'd3279015720;
		#1		read = 32'd3297210747;
		#1		read = 32'd3315290803;
		#1		read = 32'd3333254078;
		#1		read = 32'd3351098777;
		#1		read = 32'd3368823116;
		#1		read = 32'd3386425322;
		#1		read = 32'd3403903635;
		#1		read = 32'd3421256307;
		#1		read = 32'd3438481603;
		#1		read = 32'd3455577800;
		#1		read = 32'd3472543188;
		#1		read = 32'd3489376072;
		#1		read = 32'd3506074768;
		#1		read = 32'd3522637605;
		#1		read = 32'd3539062929;
		#1		read = 32'd3555349095;
		#1		read = 32'd3571494476;
		#1		read = 32'd3587497458;
		#1		read = 32'd3603356439;
		#1		read = 32'd3619069834;
		#1		read = 32'd3634636072;
		#1		read = 32'd3650053596;
		#1		read = 32'd3665320864;
		#1		read = 32'd3680436349;
		#1		read = 32'd3695398541;
		#1		read = 32'd3710205942;
		#1		read = 32'd3724857072;
		#1		read = 32'd3739350467;
		#1		read = 32'd3753684676;
		#1		read = 32'd3767858266;
		#1		read = 32'd3781869820;
		#1		read = 32'd3795717937;
		#1		read = 32'd3809401232;
		#1		read = 32'd3822918336;
		#1		read = 32'd3836267899;
		#1		read = 32'd3849448584;
		#1		read = 32'd3862459075;
		#1		read = 32'd3875298069;
		#1		read = 32'd3887964283;
		#1		read = 32'd3900456450;
		#1		read = 32'd3912773322;
		#1		read = 32'd3924913666;
		#1		read = 32'd3936876269;
		#1		read = 32'd3948659934;
		#1		read = 32'd3960263483;
		#1		read = 32'd3971685755;
		#1		read = 32'd3982925609;
		#1		read = 32'd3993981920;
		#1		read = 32'd4004853583;
		#1		read = 32'd4015539510;
		#1		read = 32'd4026038633;
		#1		read = 32'd4036349903;
		#1		read = 32'd4046472287;
		#1		read = 32'd4056404774;
		#1		read = 32'd4066146370;
		#1		read = 32'd4075696102;
		#1		read = 32'd4085053014;
		#1		read = 32'd4094216171;
		#1		read = 32'd4103184656;
		#1		read = 32'd4111957573;
		#1		read = 32'd4120534044;
		#1		read = 32'd4128913211;
		#1		read = 32'd4137094238;
		#1		read = 32'd4145076305;
		#1		read = 32'd4152858614;
		#1		read = 32'd4160440387;
		#1		read = 32'd4167820867;
		#1		read = 32'd4174999314;
		#1		read = 32'd4181975012;
		#1		read = 32'd4188747262;
		#1		read = 32'd4195315387;
		#1		read = 32'd4201678731;
		#1		read = 32'd4207836657;
		#1		read = 32'd4213788550;
		#1		read = 32'd4219533814;
		#1		read = 32'd4225071874;
		#1		read = 32'd4230402178;
		#1		read = 32'd4235524191;
		#1		read = 32'd4240437402;
		#1		read = 32'd4245141319;
		#1		read = 32'd4249635473;
		#1		read = 32'd4253919413;
		#1		read = 32'd4257992711;
		#1		read = 32'd4261854960;
		#1		read = 32'd4265505773;
		#1		read = 32'd4268944786;
		#1		read = 32'd4272171655;
		#1		read = 32'd4275186057;
		#1		read = 32'd4277987690;
		#1		read = 32'd4280576275;
		#1		read = 32'd4282951552;
		#1		read = 32'd4285113284;
		#1		read = 32'd4287061255;
		#1		read = 32'd4288795270;
		#1		read = 32'd4290315156;
		#1		read = 32'd4291620760;
		#1		read = 32'd4292711952;
		#1		read = 32'd4293588624;
		#1		read = 32'd4294250686;
		#1		read = 32'd4294698074;
		#1		read = 32'd4294930742;
		#1		read = 32'd4294948667;
		#1		read = 32'd4294751847;
		#1		read = 32'd4294340303;
		#1		read = 32'd4293714074;
		#1		read = 32'd4292873224;
		#1		read = 32'd4291817837;
		#1		read = 32'd4290548019;
		#1		read = 32'd4289063896;
		#1		read = 32'd4287365616;
		#1		read = 32'd4285453350;
		#1		read = 32'd4283327289;
		#1		read = 32'd4280987646;
		#1		read = 32'd4278434653;
		#1		read = 32'd4275668568;
		#1		read = 32'd4272689665;
		#1		read = 32'd4269498244;
		#1		read = 32'd4266094623;
		#1		read = 32'd4262479143;
		#1		read = 32'd4258652165;
		#1		read = 32'd4254614072;
		#1		read = 32'd4250365268;
		#1		read = 32'd4245906177;
		#1		read = 32'd4241237246;
		#1		read = 32'd4236358941;
		#1		read = 32'd4231271750;
		#1		read = 32'd4225976182;
		#1		read = 32'd4220472767;
		#1		read = 32'd4214762055;
		#1		read = 32'd4208844616;
		#1		read = 32'd4202721043;
		#1		read = 32'd4196391948;
		#1		read = 32'd4189857964;
		#1		read = 32'd4183119744;
		#1		read = 32'd4176177963;
		#1		read = 32'd4169033313;
		#1		read = 32'd4161686510;
		#1		read = 32'd4154138289;
		#1		read = 32'd4146389404;
		#1		read = 32'd4138440630;
		#1		read = 32'd4130292762;
		#1		read = 32'd4121946614;
		#1		read = 32'd4113403022;
		#1		read = 32'd4104662840;
		#1		read = 32'd4095726941;
		#1		read = 32'd4086596220;
		#1		read = 32'd4077271589;
		#1		read = 32'd4067753981;
		#1		read = 32'd4058044348;
		#1		read = 32'd4048143659;
		#1		read = 32'd4038052907;
		#1		read = 32'd4027773099;
		#1		read = 32'd4017305264;
		#1		read = 32'd4006650448;
		#1		read = 32'd3995809717;
		#1		read = 32'd3984784155;
		#1		read = 32'd3973574865;
		#1		read = 32'd3962182967;
		#1		read = 32'd3950609600;
		#1		read = 32'd3938855923;
		#1		read = 32'd3926923109;
		#1		read = 32'd3914812353;
		#1		read = 32'd3902524866;
		#1		read = 32'd3890061876;
		#1		read = 32'd3877424630;
		#1		read = 32'd3864614391;
		#1		read = 32'd3851632441;
		#1		read = 32'd3838480077;
		#1		read = 32'd3825158614;
		#1		read = 32'd3811669386;
		#1		read = 32'd3798013740;
		#1		read = 32'd3784193043;
		#1		read = 32'd3770208677;
		#1		read = 32'd3756062039;
		#1		read = 32'd3741754544;
		#1		read = 32'd3727287624;
		#1		read = 32'd3712662725;
		#1		read = 32'd3697881309;
		#1		read = 32'd3682944855;
		#1		read = 32'd3667854856;
		#1		read = 32'd3652612821;
		#1		read = 32'd3637220274;
		#1		read = 32'd3621678755;
		#1		read = 32'd3605989818;
		#1		read = 32'd3590155031;
		#1		read = 32'd3574175978;
		#1		read = 32'd3558054257;
		#1		read = 32'd3541791481;
		#1		read = 32'd3525389274;
		#1		read = 32'd3508849279;
		#1		read = 32'd3492173148;
		#1		read = 32'd3475362549;
		#1		read = 32'd3458419163;
		#1		read = 32'd3441344685;
		#1		read = 32'd3424140822;
		#1		read = 32'd3406809294;
		#1		read = 32'd3389351834;
		#1		read = 32'd3371770189;
		#1		read = 32'd3354066116;
		#1		read = 32'd3336241386;
		#1		read = 32'd3318297782;
		#1		read = 32'd3300237096;
		#1		read = 32'd3282061137;
		#1		read = 32'd3263771720;
		#1		read = 32'd3245370676;
		#1		read = 32'd3226859844;
		#1		read = 32'd3208241075;
		#1		read = 32'd3189516231;
		#1		read = 32'd3170687185;
		#1		read = 32'd3151755820;
		#1		read = 32'd3132724028;
		#1		read = 32'd3113593713;
		#1		read = 32'd3094366787;
		#1		read = 32'd3075045174;
		#1		read = 32'd3055630806;
		#1		read = 32'd3036125624;
		#1		read = 32'd3016531578;
		#1		read = 32'd2996850629;
		#1		read = 32'd2977084743;
		#1		read = 32'd2957235898;
		#1		read = 32'd2937306078;
		#1		read = 32'd2917297277;
		#1		read = 32'd2897211495;
		#1		read = 32'd2877050740;
		#1		read = 32'd2856817030;
		#1		read = 32'd2836512387;
		#1		read = 32'd2816138842;
		#1		read = 32'd2795698431;
		#1		read = 32'd2775193200;
		#1		read = 32'd2754625199;
		#1		read = 32'd2733996483;
		#1		read = 32'd2713309117;
		#1		read = 32'd2692565169;
		#1		read = 32'd2671766713;
		#1		read = 32'd2650915829;
		#1		read = 32'd2630014603;
		#1		read = 32'd2609065124;
		#1		read = 32'd2588069487;
		#1		read = 32'd2567029791;
		#1		read = 32'd2545948142;
		#1		read = 32'd2524826646;
		#1		read = 32'd2503667417;
		#1		read = 32'd2482472569;
		#1		read = 32'd2461244223;
		#1		read = 32'd2439984501;
		#1		read = 32'd2418695529;
		#1		read = 32'd2397379436;
		#1		read = 32'd2376038354;
		#1		read = 32'd2354674416;
		#1		read = 32'd2333289760;
		#1		read = 32'd2311886523;
		#1		read = 32'd2290466846;
		#1		read = 32'd2269032871;
		#1		read = 32'd2247586740;
		#1		read = 32'd2226130600;
		#1		read = 32'd2204666595;
		#1		read = 32'd2183196872;
		#1		read = 32'd2161723578;
		#1		read = 32'd2140248859;
		#1		read = 32'd2118774864;
		#1		read = 32'd2097303740;
		#1		read = 32'd2075837634;
		#1		read = 32'd2054378692;
		#1		read = 32'd2032929061;
		#1		read = 32'd2011490885;
		#1		read = 32'd1990066309;
		#1		read = 32'd1968657474;
		#1		read = 32'd1947266521;
		#1		read = 32'd1925895590;
		#1		read = 32'd1904546817;
		#1		read = 32'd1883222339;
		#1		read = 32'd1861924285;
		#1		read = 32'd1840654788;
		#1		read = 32'd1819415973;
		#1		read = 32'd1798209965;
		#1		read = 32'd1777038884;
		#1		read = 32'd1755904847;
		#1		read = 32'd1734809968;
		#1		read = 32'd1713756355;
		#1		read = 32'd1692746115;
		#1		read = 32'd1671781349;
		#1		read = 32'd1650864152;
		#1		read = 32'd1629996616;
		#1		read = 32'd1609180829;
		#1		read = 32'd1588418872;
		#1		read = 32'd1567712821;
		#1		read = 32'd1547064746;
		#1		read = 32'd1526476713;
		#1		read = 32'd1505950780;
		#1		read = 32'd1485489000;
		#1		read = 32'd1465093419;
		#1		read = 32'd1444766076;
		#1		read = 32'd1424509004;
		#1		read = 32'd1404324229;
		#1		read = 32'd1384213770;
		#1		read = 32'd1364179637;
		#1		read = 32'd1344223833;
		#1		read = 32'd1324348355;
		#1		read = 32'd1304555190;
		#1		read = 32'd1284846317;
		#1		read = 32'd1265223706;
		#1		read = 32'd1245689322;
		#1		read = 32'd1226245115;
		#1		read = 32'd1206893032;
		#1		read = 32'd1187635008;
		#1		read = 32'd1168472967;
		#1		read = 32'd1149408826;
		#1		read = 32'd1130444492;
		#1		read = 32'd1111581862;
		#1		read = 32'd1092822820;
		#1		read = 32'd1074169244;
		#1		read = 32'd1055622998;
		#1		read = 32'd1037185938;
		#1		read = 32'd1018859906;
		#1		read = 32'd1000646736;
		#1		read = 32'd982548248;
		#1		read = 32'd964566253;
		#1		read = 32'd946702549;
		#1		read = 32'd928958922;
		#1		read = 32'd911337146;
		#1		read = 32'd893838984;
		#1		read = 32'd876466185;
		#1		read = 32'd859220488;
		#1		read = 32'd842103615;
		#1		read = 32'd825117279;
		#1		read = 32'd808263179;
		#1		read = 32'd791543000;
		#1		read = 32'd774958413;
		#1		read = 32'd758511078;
		#1		read = 32'd742202639;
		#1		read = 32'd726034727;
		#1		read = 32'd710008959;
		#1		read = 32'd694126937;
		#1		read = 32'd678390250;
		#1		read = 32'd662800470;
		#1		read = 32'd647359158;
		#1		read = 32'd632067857;
		#1		read = 32'd616928096;
		#1		read = 32'd601941389;
		#1		read = 32'd587109236;
		#1		read = 32'd572433118;
		#1		read = 32'd557914505;
		#1		read = 32'd543554847;
		#1		read = 32'd529355580;
		#1		read = 32'd515318125;
		#1		read = 32'd501443885;
		#1		read = 32'd487734248;
		#1		read = 32'd474190584;
		#1		read = 32'd460814248;
		#1		read = 32'd447606578;
		#1		read = 32'd434568894;
		#1		read = 32'd421702500;
		#1		read = 32'd409008682;
		#1		read = 32'd396488711;
		#1		read = 32'd384143838;
		#1		read = 32'd371975297;
		#1		read = 32'd359984306;
		#1		read = 32'd348172063;
		#1		read = 32'd336539750;
		#1		read = 32'd325088529;
		#1		read = 32'd313819547;
		#1		read = 32'd302733929;
		#1		read = 32'd291832785;
		#1		read = 32'd281117205;
		#1		read = 32'd270588259;
		#1		read = 32'd260247002;
		#1		read = 32'd250094467;
		#1		read = 32'd240131669;
		#1		read = 32'd230359604;
		#1		read = 32'd220779251;
		#1		read = 32'd211391566;
		#1		read = 32'd202197489;
		#1		read = 32'd193197938;
		#1		read = 32'd184393815;
		#1		read = 32'd175785999;
		#1		read = 32'd167375352;
		#1		read = 32'd159162713;
		#1		read = 32'd151148905;
		#1		read = 32'd143334728;
		#1		read = 32'd135720965;
		#1		read = 32'd128308377;
		#1		read = 32'd121097704;
		#1		read = 32'd114089668;
		#1		read = 32'd107284970;
		#1		read = 32'd100684290;
		#1		read = 32'd94288289;
		#1		read = 32'd88097605;
		#1		read = 32'd82112858;
		#1		read = 32'd76334646;
		#1		read = 32'd70763548;
		#1		read = 32'd65400120;
		#1		read = 32'd60244898;
		#1		read = 32'd55298399;
		#1		read = 32'd50561116;
		#1		read = 32'd46033524;
		#1		read = 32'd41716075;
		#1		read = 32'd37609201;
		#1		read = 32'd33713313;
		#1		read = 32'd30028800;
		#1		read = 32'd26556031;
		#1		read = 32'd23295353;
		#1		read = 32'd20247092;
		#1		read = 32'd17411552;
		#1		read = 32'd14789019;
		#1		read = 32'd12379752;
		#1		read = 32'd10183995;
		#1		read = 32'd8201966;
		#1		read = 32'd6433863;
		#1		read = 32'd4879863;
		#1		read = 32'd3540122;
		#1		read = 32'd2414773;
		#1		read = 32'd1503930;
		#1		read = 32'd807682;
		#1		read = 32'd326101;
		#1		read = 32'd59233;
		#1		read = 32'd7107;
		#1		read = 32'd169726;
		#1		read = 32'd547074;
		#1		read = 32'd1139115;
		#1		read = 32'd1945788;
		#1		read = 32'd2967013;
		#1		read = 32'd4202688;
		#1		read = 32'd5652689;
		#1		read = 32'd7316872;
		#1		read = 32'd9195069;
		#1		read = 32'd11287094;
		#1		read = 32'd13592736;
		#1		read = 32'd16111766;
		#1		read = 32'd18843931;
		#1		read = 32'd21788959;
		#1		read = 32'd24946554;
		#1		read = 32'd28316401;
		#1		read = 32'd31898163;
		#1		read = 32'd35691482;
		#1		read = 32'd39695978;
		#1		read = 32'd43911251;
		#1		read = 32'd48336880;
		#1		read = 32'd52972421;
		#1		read = 32'd57817412;
		#1		read = 32'd62871368;
		#1		read = 32'd68133784;
		#1		read = 32'd73604132;
		#1		read = 32'd79281867;
		#1		read = 32'd85166421;
		#1		read = 32'd91257204;
		#1		read = 32'd97553608;
		#1		read = 32'd104055004;
		#1		read = 32'd110760740;
		#1		read = 32'd117670148;
		#1		read = 32'd124782535;
		#1		read = 32'd132097190;
		#1		read = 32'd139613383;
		#1		read = 32'd147330360;
		#1		read = 32'd155247352;
		#1		read = 32'd163363565;
		#1		read = 32'd171678189;
		#1		read = 32'd180190391;
		#1		read = 32'd188899322;
		#1		read = 32'd197804109;
		#1		read = 32'd206903862;
		#1		read = 32'd216197672;
		#1		read = 32'd225684609;
		#1		read = 32'd235363724;
		#1		read = 32'd245234049;
		#1		read = 32'd255294598;
		#1		read = 32'd265544364;
		#1		read = 32'd275982323;
		#1		read = 32'd286607430;
		#1		read = 32'd297418623;
		#1		read = 32'd308414821;
		#1		read = 32'd319594925;
		#1		read = 32'd330957816;
		#1		read = 32'd342502357;
		#1		read = 32'd354227396;
		#1		read = 32'd366131759;
		#1		read = 32'd378214255;
		#1		read = 32'd390473677;
		#1		read = 32'd402908798;
		#1		read = 32'd415518376;
		#1		read = 32'd428301148;
		#1		read = 32'd441255837;
		#1		read = 32'd454381148;
		#1		read = 32'd467675768;
		#1		read = 32'd481138367;
		#1		read = 32'd494767599;
		#1		read = 32'd508562101;
		#1		read = 32'd522520494;
		#1		read = 32'd536641382;
		#1		read = 32'd550923353;
		#1		read = 32'd565364978;
		#1		read = 32'd579964814;
		#1		read = 32'd594721401;
		#1		read = 32'd609633263;
		#1		read = 32'd624698908;
		#1		read = 32'd639916831;
		#1		read = 32'd655285509;
		#1		read = 32'd670803405;
		#1		read = 32'd686468969;
		#1		read = 32'd702280633;
		#1		read = 32'd718236815;
		#1		read = 32'd734335922;
		#1		read = 32'd750576341;
		#1		read = 32'd766956451;
		#1		read = 32'd783474612;
		#1		read = 32'd800129172;
		#1		read = 32'd816918468;
		#1		read = 32'd833840818;
		#1		read = 32'd850894532;
		#1		read = 32'd868077903;
		#1		read = 32'd885389214;
		#1		read = 32'd902826734;
		#1		read = 32'd920388718;
		#1		read = 32'd938073410;
		#1		read = 32'd955879043;
		#1		read = 32'd973803835;
		#1		read = 32'd991845994;
		#1		read = 32'd1010003715;
		#1		read = 32'd1028275184;
		#1		read = 32'd1046658573;
		#1		read = 32'd1065152043;
		#1		read = 32'd1083753746;
		#1		read = 32'd1102461821;
		#1		read = 32'd1121274397;
		#1		read = 32'd1140189593;
		#1		read = 32'd1159205517;
		#1		read = 32'd1178320269;
		#1		read = 32'd1197531936;
		#1		read = 32'd1216838598;
		#1		read = 32'd1236238323;
		#1		read = 32'd1255729172;
		#1		read = 32'd1275309196;
		#1		read = 32'd1294976436;
		#1		read = 32'd1314728927;
		#1		read = 32'd1334564692;
		#1		read = 32'd1354481749;
		#1		read = 32'd1374478105;
		#1		read = 32'd1394551761;
		#1		read = 32'd1414700709;
		#1		read = 32'd1434922935;
		#1		read = 32'd1455216417;
		#1		read = 32'd1475579125;
		#1		read = 32'd1496009023;
		#1		read = 32'd1516504067;
		#1		read = 32'd1537062209;
		#1		read = 32'd1557681393;
		#1		read = 32'd1578359556;
		#1		read = 32'd1599094632;
		#1		read = 32'd1619884545;
		#1		read = 32'd1640727219;
		#1		read = 32'd1661620567;
		#1		read = 32'd1682562502;
		#1		read = 32'd1703550928;
		#1		read = 32'd1724583747;
		#1		read = 32'd1745658855;
		#1		read = 32'd1766774146;
		#1		read = 32'd1787927508;
		#1		read = 32'd1809116824;
		#1		read = 32'd1830339977;
		#1		read = 32'd1851594845;
		#1		read = 32'd1872879301;
		#1		read = 32'd1894191217;
		#1		read = 32'd1915528462;
		#1		read = 32'd1936888902;
		#1		read = 32'd1958270402;
		#1		read = 32'd1979670823;
		#1		read = 32'd2001088025;
		#1		read = 32'd2022519866;
		#1		read = 32'd2043964204;
		#1		read = 32'd2065418894;
		#1		read = 32'd2086881790;
		#1		read = 32'd2108350746;
		#1		read = 32'd2129823616;
		#1		read = 32'd2151298251;
		#1		read = 32'd2172772505;
		#1		read = 32'd2194244230;
		#1		read = 32'd2215711279;
		#1		read = 32'd2237171505;
		#1		read = 32'd2258622763;
		#1		read = 32'd2280062907;
		#1		read = 32'd2301489793;
		#1		read = 32'd2322901278;
		#1		read = 32'd2344295222;
		#1		read = 32'd2365669485;
		#1		read = 32'd2387021930;
		#1		read = 32'd2408350421;
		#1		read = 32'd2429652825;
		#1		read = 32'd2450927013;
		#1		read = 32'd2472170857;
		#1		read = 32'd2493382232;
		#1		read = 32'd2514559018;
		#1		read = 32'd2535699096;
		#1		read = 32'd2556800353;
		#1		read = 32'd2577860679;
		#1		read = 32'd2598877968;
		#1		read = 32'd2619850117;
		#1		read = 32'd2640775030;
		#1		read = 32'd2661650615;
		#1		read = 32'd2682474783;
		#1		read = 32'd2703245452;
		#1		read = 32'd2723960546;
		#1		read = 32'd2744617993;
		#1		read = 32'd2765215727;
		#1		read = 32'd2785751688;
		#1		read = 32'd2806223822;
		#1		read = 32'd2826630084;
		#1		read = 32'd2846968431;
		#1		read = 32'd2867236830;
		#1		read = 32'd2887433255;
		#1		read = 32'd2907555685;
		#1		read = 32'd2927602108;
		#1		read = 32'd2947570521;
		#1		read = 32'd2967458925;
		#1		read = 32'd2987265333;
		#1		read = 32'd3006987763;
		#1		read = 32'd3026624244;
		#1		read = 32'd3046172811;
		#1		read = 32'd3065631510;
		#1		read = 32'd3084998394;
		#1		read = 32'd3104271529;
		#1		read = 32'd3123448985;
		#1		read = 32'd3142528845;
		#1		read = 32'd3161509202;
		#1		read = 32'd3180388157;
		#1		read = 32'd3199163823;
		#1		read = 32'd3217834321;
		#1		read = 32'd3236397785;
		#1		read = 32'd3254852359;
		#1		read = 32'd3273196197;
		#1		read = 32'd3291427464;
		#1		read = 32'd3309544338;
		#1		read = 32'd3327545007;
		#1		read = 32'd3345427671;
		#1		read = 32'd3363190541;
		#1		read = 32'd3380831842;
		#1		read = 32'd3398349809;
		#1		read = 32'd3415742690;
		#1		read = 32'd3433008747;
		#1		read = 32'd3450146252;
		#1		read = 32'd3467153491;
		#1		read = 32'd3484028765;
		#1		read = 32'd3500770386;
		#1		read = 32'd3517376679;
		#1		read = 32'd3533845984;
		#1		read = 32'd3550176654;
		#1		read = 32'd3566367055;
		#1		read = 32'd3582415570;
		#1		read = 32'd3598320592;
		#1		read = 32'd3614080532;
		#1		read = 32'd3629693814;
		#1		read = 32'd3645158875;
		#1		read = 32'd3660474171;
		#1		read = 32'd3675638169;
		#1		read = 32'd3690649352;
		#1		read = 32'd3705506220;
		#1		read = 32'd3720207288;
		#1		read = 32'd3734751084;
		#1		read = 32'd3749136155;
		#1		read = 32'd3763361061;
		#1		read = 32'd3777424382;
		#1		read = 32'd3791324710;
		#1		read = 32'd3805060655;
		#1		read = 32'd3818630843;
		#1		read = 32'd3832033919;
		#1		read = 32'd3845268541;
		#1		read = 32'd3858333385;
		#1		read = 32'd3871227146;
		#1		read = 32'd3883948535;
		#1		read = 32'd3896496278;
		#1		read = 32'd3908869121;
		#1		read = 32'd3921065827;
		#1		read = 32'd3933085177;
		#1		read = 32'd3944925968;
		#1		read = 32'd3956587016;
		#1		read = 32'd3968067155;
		#1		read = 32'd3979365238;
		#1		read = 32'd3990480134;
		#1		read = 32'd4001410731;
		#1		read = 32'd4012155938;
		#1		read = 32'd4022714679;
		#1		read = 32'd4033085898;
		#1		read = 32'd4043268559;
		#1		read = 32'd4053261643;
		#1		read = 32'd4063064150;
		#1		read = 32'd4072675102;
		#1		read = 32'd4082093535;
		#1		read = 32'd4091318509;
		#1		read = 32'd4100349102;
		#1		read = 32'd4109184409;
		#1		read = 32'd4117823548;
		#1		read = 32'd4126265655;
		#1		read = 32'd4134509885;
		#1		read = 32'd4142555414;
		#1		read = 32'd4150401438;
		#1		read = 32'd4158047171;
		#1		read = 32'd4165491850;
		#1		read = 32'd4172734730;
		#1		read = 32'd4179775086;
		#1		read = 32'd4186612215;
		#1		read = 32'd4193245432;
		#1		read = 32'd4199674076;
		#1		read = 32'd4205897501;
		#1		read = 32'd4211915088;
		#1		read = 32'd4217726232;
		#1		read = 32'd4223330355;
		#1		read = 32'd4228726894;
		#1		read = 32'd4233915311;
		#1		read = 32'd4238895086;
		#1		read = 32'd4243665722;
		#1		read = 32'd4248226741;
		#1		read = 32'd4252577688;
		#1		read = 32'd4256718127;
		#1		read = 32'd4260647645;
		#1		read = 32'd4264365848;
		#1		read = 32'd4267872364;
		#1		read = 32'd4271166843;
		#1		read = 32'd4274248956;
		#1		read = 32'd4277118394;
		#1		read = 32'd4279774870;
		#1		read = 32'd4282218119;
		#1		read = 32'd4284447897;
		#1		read = 32'd4286463979;
		#1		read = 32'd4288266166;
		#1		read = 32'd4289854276;
		#1		read = 32'd4291228150;
		#1		read = 32'd4292387652;
		#1		read = 32'd4293332666;
		#1		read = 32'd4294063096;
		#1		read = 32'd4294578870;
		#1		read = 32'd4294879936;
		#1		read = 32'd4294966265;
		#1		read = 32'd4294837847;
		#1		read = 32'd4294494695;
		#1		read = 32'd4293936844;
		#1		read = 32'd4293164350;
		#1		read = 32'd4292177289;
		#1		read = 32'd4290975761;
		#1		read = 32'd4289559885;
		#1		read = 32'd4287929804;
		#1		read = 32'd4286085679;
		#1		read = 32'd4284027697;
		#1		read = 32'd4281756061;
		#1		read = 32'd4279271000;
		#1		read = 32'd4276572762;
		#1		read = 32'd4273661617;
		#1		read = 32'd4270537856;
		#1		read = 32'd4267201792;
		#1		read = 32'd4263653757;
		#1		read = 32'd4259894107;
		#1		read = 32'd4255923218;
		#1		read = 32'd4251741486;
		#1		read = 32'd4247349331;
		#1		read = 32'd4242747191;
		#1		read = 32'd4237935526;
		#1		read = 32'd4232914817;
		#1		read = 32'd4227685568;
		#1		read = 32'd4222248300;
		#1		read = 32'd4216603557;
		#1		read = 32'd4210751903;
		#1		read = 32'd4204693925;
		#1		read = 32'd4198430228;
		#1		read = 32'd4191961437;
		#1		read = 32'd4185288200;
		#1		read = 32'd4178411185;
		#1		read = 32'd4171331079;
		#1		read = 32'd4164048589;
		#1		read = 32'd4156564445;
		#1		read = 32'd4148879394;
		#1		read = 32'd4140994205;
		#1		read = 32'd4132909667;
		#1		read = 32'd4124626588;
		#1		read = 32'd4116145797;
		#1		read = 32'd4107468141;
		#1		read = 32'd4098594488;
		#1		read = 32'd4089525725;
		#1		read = 32'd4080262760;
		#1		read = 32'd4070806519;
		#1		read = 32'd4061157947;
		#1		read = 32'd4051318009;
		#1		read = 32'd4041287689;
		#1		read = 32'd4031067991;
		#1		read = 32'd4020659935;
		#1		read = 32'd4010064564;
		#1		read = 32'd3999282936;
		#1		read = 32'd3988316129;
		#1		read = 32'd3977165241;
		#1		read = 32'd3965831386;
		#1		read = 32'd3954315698;
		#1		read = 32'd3942619329;
		#1		read = 32'd3930743447;
		#1		read = 32'd3918689241;
		#1		read = 32'd3906457915;
		#1		read = 32'd3894050694;
		#1		read = 32'd3881468817;
		#1		read = 32'd3868713544;
		#1		read = 32'd3855786149;
		#1		read = 32'd3842687925;
		#1		read = 32'd3829420182;
		#1		read = 32'd3815984246;
		#1		read = 32'd3802381462;
		#1		read = 32'd3788613190;
		#1		read = 32'd3774680806;
		#1		read = 32'd3760585704;
		#1		read = 32'd3746329292;
		#1		read = 32'd3731912998;
		#1		read = 32'd3717338262;
		#1		read = 32'd3702606542;
		#1		read = 32'd3687719311;
		#1		read = 32'd3672678057;
		#1		read = 32'd3657484286;
		#1		read = 32'd3642139515;
		#1		read = 32'd3626645280;
		#1		read = 32'd3611003131;
		#1		read = 32'd3595214630;
		#1		read = 32'd3579281358;
		#1		read = 32'd3563204907;
		#1		read = 32'd3546986885;
		#1		read = 32'd3530628914;
		#1		read = 32'd3514132630;
		#1		read = 32'd3497499682;
		#1		read = 32'd3480731733;
		#1		read = 32'd3463830461;
		#1		read = 32'd3446797555;
		#1		read = 32'd3429634719;
		#1		read = 32'd3412343669;
		#1		read = 32'd3394926133;
		#1		read = 32'd3377383855;
		#1		read = 32'd3359718588;
		#1		read = 32'd3341932098;
		#1		read = 32'd3324026164;
		#1		read = 32'd3306002577;
		#1		read = 32'd3287863139;
		#1		read = 32'd3269609664;
		#1		read = 32'd3251243978;
		#1		read = 32'd3232767916;
		#1		read = 32'd3214183327;
		#1		read = 32'd3195492068;
		#1		read = 32'd3176696010;
		#1		read = 32'd3157797032;
		#1		read = 32'd3138797022;
		#1		read = 32'd3119697883;
		#1		read = 32'd3100501522;
		#1		read = 32'd3081209861;
		#1		read = 32'd3061824828;
		#1		read = 32'd3042348362;
		#1		read = 32'd3022782409;
		#1		read = 32'd3003128928;
		#1		read = 32'd2983389883;
		#1		read = 32'd2963567248;
		#1		read = 32'd2943663005;
		#1		read = 32'd2923679145;
		#1		read = 32'd2903617666;
		#1		read = 32'd2883480574;
		#1		read = 32'd2863269884;
		#1		read = 32'd2842987615;
		#1		read = 32'd2822635796;
		#1		read = 32'd2802216463;
		#1		read = 32'd2781731657;
		#1		read = 32'd2761183427;
		#1		read = 32'd2740573827;
		#1		read = 32'd2719904919;
		#1		read = 32'd2699178769;
		#1		read = 32'd2678397450;
		#1		read = 32'd2657563040;
		#1		read = 32'd2636677622;
		#1		read = 32'd2615743286;
		#1		read = 32'd2594762124;
		#1		read = 32'd2573736235;
		#1		read = 32'd2552667720;
		#1		read = 32'd2531558688;
		#1		read = 32'd2510411248;
		#1		read = 32'd2489227516;
		#1		read = 32'd2468009610;
		#1		read = 32'd2446759651;
		#1		read = 32'd2425479765;
		#1		read = 32'd2404172080;
		#1		read = 32'd2382838726;
		#1		read = 32'd2361481837;
		#1		read = 32'd2340103548;
		#1		read = 32'd2318705998;
		#1		read = 32'd2297291325;
		#1		read = 32'd2275861672;
		#1		read = 32'd2254419180;
		#1		read = 32'd2232965996;
		#1		read = 32'd2211504263;
		#1		read = 32'd2190036128;
		#1		read = 32'd2168563739;
		#1		read = 32'd2147089241;
		#1		read = 32'd2125614782;
		#1		read = 32'd2104142511;
		#1		read = 32'd2082674573;
		#1		read = 32'd2061213116;
		#1		read = 32'd2039760287;
		#1		read = 32'd2018318229;
		#1		read = 32'd1996889088;
		#1		read = 32'd1975475006;
		#1		read = 32'd1954078125;
		#1		read = 32'd1932700585;
		#1		read = 32'd1911344522;
		#1		read = 32'd1890012074;
		#1		read = 32'd1868705372;
		#1		read = 32'd1847426548;
		#1		read = 32'd1826177729;
		#1		read = 32'd1804961040;
		#1		read = 32'd1783778604;
		#1		read = 32'd1762632538;
		#1		read = 32'd1741524956;
		#1		read = 32'd1720457970;
		#1		read = 32'd1699433687;
		#1		read = 32'd1678454208;
		#1		read = 32'd1657521631;
		#1		read = 32'd1636638050;
		#1		read = 32'd1615805554;
		#1		read = 32'd1595026225;
		#1		read = 32'd1574302141;
		#1		read = 32'd1553635374;
		#1		read = 32'd1533027992;
		#1		read = 32'd1512482055;
		#1		read = 32'd1491999618;
		#1		read = 32'd1471582729;
		#1		read = 32'd1451233429;
		#1		read = 32'd1430953753;
		#1		read = 32'd1410745730;
		#1		read = 32'd1390611381;
		#1		read = 32'd1370552717;
		#1		read = 32'd1350571746;
		#1		read = 32'd1330670466;
		#1		read = 32'd1310850867;
		#1		read = 32'd1291114929;
		#1		read = 32'd1271464628;
		#1		read = 32'd1251901929;
		#1		read = 32'd1232428786;
		#1		read = 32'd1213047149;
		#1		read = 32'd1193758954;
		#1		read = 32'd1174566131;
		#1		read = 32'd1155470599;
		#1		read = 32'd1136474267;
		#1		read = 32'd1117579036;
		#1		read = 32'd1098786794;
		#1		read = 32'd1080099421;
		#1		read = 32'd1061518785;
		#1		read = 32'd1043046745;
		#1		read = 32'd1024685148;
		#1		read = 32'd1006435829;
		#1		read = 32'd988300615;
		#1		read = 32'd970281318;
		#1		read = 32'd952379740;
		#1		read = 32'd934597671;
		#1		read = 32'd916936890;
		#1		read = 32'd899399163;
		#1		read = 32'd881986243;
		#1		read = 32'd864699872;
		#1		read = 32'd847541778;
		#1		read = 32'd830513678;
		#1		read = 32'd813617273;
		#1		read = 32'd796854253;
		#1		read = 32'd780226296;
		#1		read = 32'd763735063;
		#1		read = 32'd747382204;
		#1		read = 32'd731169353;
		#1		read = 32'd715098133;
		#1		read = 32'd699170151;
		#1		read = 32'd683386998;
		#1		read = 32'd667750254;
		#1		read = 32'd652261482;
		#1		read = 32'd636922231;
		#1		read = 32'd621734035;
		#1		read = 32'd606698413;
		#1		read = 32'd591816868;
		#1		read = 32'd577090888;
		#1		read = 32'd562521946;
		#1		read = 32'd548111499;
		#1		read = 32'd533860988;
		#1		read = 32'd519771838;
		#1		read = 32'd505845457;
		#1		read = 32'd492083239;
		#1		read = 32'd478486560;
		#1		read = 32'd465056779;
		#1		read = 32'd451795240;
		#1		read = 32'd438703268;
		#1		read = 32'd425782172;
		#1		read = 32'd413033245;
		#1		read = 32'd400457762;
		#1		read = 32'd388056980;
		#1		read = 32'd375832139;
		#1		read = 32'd363784461;
		#1		read = 32'd351915153;
		#1		read = 32'd340225399;
		#1		read = 32'd328716370;
		#1		read = 32'd317389216;
		#1		read = 32'd306245070;
		#1		read = 32'd295285046;
		#1		read = 32'd284510241;
		#1		read = 32'd273921731;
		#1		read = 32'd263520576;
		#1		read = 32'd253307816;
		#1		read = 32'd243284472;
		#1		read = 32'd233451546;
		#1		read = 32'd223810022;
		#1		read = 32'd214360863;
		#1		read = 32'd205105015;
		#1		read = 32'd196043404;
		#1		read = 32'd187176934;
		#1		read = 32'd178506494;
		#1		read = 32'd170032950;
		#1		read = 32'd161757149;
		#1		read = 32'd153679920;
		#1		read = 32'd145802069;
		#1		read = 32'd138124384;
		#1		read = 32'd130647634;
		#1		read = 32'd123372566;
		#1		read = 32'd116299907;
		#1		read = 32'd109430365;
		#1		read = 32'd102764626;
		#1		read = 32'd96303358;
		#1		read = 32'd90047206;
		#1		read = 32'd83996795;
		#1		read = 32'd78152732;
		#1		read = 32'd72515601;
		#1		read = 32'd67085964;
		#1		read = 32'd61864365;
		#1		read = 32'd56851327;
		#1		read = 32'd52047350;
		#1		read = 32'd47452914;
		#1		read = 32'd43068481;
		#1		read = 32'd38894487;
		#1		read = 32'd34931350;
		#1		read = 32'd31179466;
		#1		read = 32'd27639212;
		#1		read = 32'd24310939;
		#1		read = 32'd21194983;
		#1		read = 32'd18291653;
		#1		read = 32'd15601241;
		#1		read = 32'd13124016;
		#1		read = 32'd10860224;
		#1		read = 32'd8810094;
		#1		read = 32'd6973828;
		#1		read = 32'd5351612;
		#1		read = 32'd3943608;
		#1		read = 32'd2749955;
		#1		read = 32'd1770774;
		#1		read = 32'd1006163;
		#1		read = 32'd456197;
		#1		read = 32'd120933;
		#1		read = 32'd403;
		#1		read = 32'd94620;
		#1		read = 32'd403573;
		#1		read = 32'd927233;
		#1		read = 32'd1665547;
		#1		read = 32'd2618441;
		#1		read = 32'd3785819;
		#1		read = 32'd5167566;
		#1		read = 32'd6763542;
		#1		read = 32'd8573589;
		#1		read = 32'd10597524;
		#1		read = 32'd12835147;
		#1		read = 32'd15286233;
		#1		read = 32'd17950536;
		#1		read = 32'd20827792;
		#1		read = 32'd23917711;
		#1		read = 32'd27219984;
		#1		read = 32'd30734283;
		#1		read = 32'd34460254;
		#1		read = 32'd38397527;
		#1		read = 32'd42545706;
		#1		read = 32'd46904377;
		#1		read = 32'd51473104;
		#1		read = 32'd56251431;
		#1		read = 32'd61238879;
		#1		read = 32'd66434949;
		#1		read = 32'd71839123;
		#1		read = 32'd77450860;
		#1		read = 32'd83269598;
		#1		read = 32'd89294756;
		#1		read = 32'd95525731;
		#1		read = 32'd101961900;
		#1		read = 32'd108602620;
		#1		read = 32'd115447226;
		#1		read = 32'd122495034;
		#1		read = 32'd129745339;
		#1		read = 32'd137197416;
		#1		read = 32'd144850520;
		#1		read = 32'd152703886;
		#1		read = 32'd160756728;
		#1		read = 32'd169008241;
		#1		read = 32'd177457601;
		#1		read = 32'd186103961;
		#1		read = 32'd194946457;
		#1		read = 32'd203984206;
		#1		read = 32'd213216302;
		#1		read = 32'd222641824;
		#1		read = 32'd232259829;
		#1		read = 32'd242069354;
		#1		read = 32'd252069419;
		#1		read = 32'd262259024;
		#1		read = 32'd272637150;
		#1		read = 32'd283202759;
		#1		read = 32'd293954795;
		#1		read = 32'd304892181;
		#1		read = 32'd316013826;
		#1		read = 32'd327318616;
		#1		read = 32'd338805421;
		#1		read = 32'd350473092;
		#1		read = 32'd362320463;
		#1		read = 32'd374346348;
		#1		read = 32'd386549546;
		#1		read = 32'd398928836;
		#1		read = 32'd411482980;
		#1		read = 32'd424210722;
		#1		read = 32'd437110791;
		#1		read = 32'd450181895;
		#1		read = 32'd463422728;
		#1		read = 32'd476831965;
		#1		read = 32'd490408267;
		#1		read = 32'd504150274;
		#1		read = 32'd518056614;
		#1		read = 32'd532125895;
		#1		read = 32'd546356710;
		#1		read = 32'd560747636;
		#1		read = 32'd575297235;
		#1		read = 32'd590004052;
		#1		read = 32'd604866615;
		#1		read = 32'd619883438;
		#1		read = 32'd635053020;
		#1		read = 32'd650373844;
		#1		read = 32'd665844377;
		#1		read = 32'd681463074;
		#1		read = 32'd697228371;
		#1		read = 32'd713138692;
		#1		read = 32'd729192447;
		#1		read = 32'd745388030;
		#1		read = 32'd761723821;
		#1		read = 32'd778198187;
		#1		read = 32'd794809480;
		#1		read = 32'd811556040;
		#1		read = 32'd828436191;
		#1		read = 32'd845448246;
		#1		read = 32'd862590503;
		#1		read = 32'd879861249;
		#1		read = 32'd897258756;
		#1		read = 32'd914781284;
		#1		read = 32'd932427081;
		#1		read = 32'd950194384;
		#1		read = 32'd968081414;
		#1		read = 32'd986086383;
		#1		read = 32'd1004207491;
		#1		read = 32'd1022442926;
		#1		read = 32'd1040790863;
		#1		read = 32'd1059249470;
		#1		read = 32'd1077816898;
		#1		read = 32'd1096491293;
		#1		read = 32'd1115270786;
		#1		read = 32'd1134153499;
		#1		read = 32'd1153137544;
		#1		read = 32'd1172221023;
		#1		read = 32'd1191402028;
		#1		read = 32'd1210678640;
		#1		read = 32'd1230048932;
		#1		read = 32'd1249510966;
		#1		read = 32'd1269062797;
		#1		read = 32'd1288702470;
		#1		read = 32'd1308428019;
		#1		read = 32'd1328237474;
		#1		read = 32'd1348128853;
		#1		read = 32'd1368100166;
		#1		read = 32'd1388149417;
		#1		read = 32'd1408274601;
		#1		read = 32'd1428473705;
		#1		read = 32'd1448744709;
		#1		read = 32'd1469085587;
		#1		read = 32'd1489494304;
		#1		read = 32'd1509968820;
		#1		read = 32'd1530507086;
		#1		read = 32'd1551107050;
		#1		read = 32'd1571766650;
		#1		read = 32'd1592483822;
		#1		read = 32'd1613256494;
		#1		read = 32'd1634082587;
		#1		read = 32'd1654960021;
		#1		read = 32'd1675886706;
		#1		read = 32'd1696860551;
		#1		read = 32'd1717879457;
		#1		read = 32'd1738941324;
		#1		read = 32'd1760044045;
		#1		read = 32'd1781185509;
		#1		read = 32'd1802363602;
		#1		read = 32'd1823576208;
		#1		read = 32'd1844821204;
		#1		read = 32'd1866096466;
		#1		read = 32'd1887399866;
		#1		read = 32'd1908729274;
		#1		read = 32'd1930082558;
		#1		read = 32'd1951457582;
		#1		read = 32'd1972852208;
		#1		read = 32'd1994264297;
		#1		read = 32'd2015691708;
		#1		read = 32'd2037132298;
		#1		read = 32'd2058583923;
		#1		read = 32'd2080044438;
		#1		read = 32'd2101511697;
		#1		read = 32'd2122983553;
		#1		read = 32'd2144457859;
		#1		read = 32'd2165932467;
		#1		read = 32'd2187405231;
		#1		read = 32'd2208874003;
		#1		read = 32'd2230336635;
		#1		read = 32'd2251790983;
		#1		read = 32'd2273234899;
		#1		read = 32'd2294666241;
		#1		read = 32'd2316082864;
		#1		read = 32'd2337482628;
		#1		read = 32'd2358863392;
		#1		read = 32'd2380223018;
		#1		read = 32'd2401559371;
		#1		read = 32'd2422870316;
		#1		read = 32'd2444153723;
		#1		read = 32'd2465407463;
		#1		read = 32'd2486629410;
		#1		read = 32'd2507817444;
		#1		read = 32'd2528969444;
		#1		read = 32'd2550083296;
		#1		read = 32'd2571156889;
		#1		read = 32'd2592188114;
		#1		read = 32'd2613174870;
		#1		read = 32'd2634115057;
		#1		read = 32'd2655006581;
		#1		read = 32'd2675847353;
		#1		read = 32'd2696635289;
		#1		read = 32'd2717368311;
		#1		read = 32'd2738044344;
		#1		read = 32'd2758661322;
		#1		read = 32'd2779217183;
		#1		read = 32'd2799709871;
		#1		read = 32'd2820137336;
		#1		read = 32'd2840497537;
		#1		read = 32'd2860788437;
		#1		read = 32'd2881008008;
		#1		read = 32'd2901154226;
		#1		read = 32'd2921225078;
		#1		read = 32'd2941218557;
		#1		read = 32'd2961132662;
		#1		read = 32'd2980965404;
		#1		read = 32'd3000714798;
		#1		read = 32'd3020378869;
		#1		read = 32'd3039955652;
		#1		read = 32'd3059443189;
		#1		read = 32'd3078839530;
		#1		read = 32'd3098142736;
		#1		read = 32'd3117350877;
		#1		read = 32'd3136462032;
		#1		read = 32'd3155474291;
		#1		read = 32'd3174385751;
		#1		read = 32'd3193194522;
		#1		read = 32'd3211898722;
		#1		read = 32'd3230496482;
		#1		read = 32'd3248985941;
		#1		read = 32'd3267365252;
		#1		read = 32'd3285632574;
		#1		read = 32'd3303786083;
		#1		read = 32'd3321823963;
		#1		read = 32'd3339744410;
		#1		read = 32'd3357545631;
		#1		read = 32'd3375225848;
		#1		read = 32'd3392783291;
		#1		read = 32'd3410216205;
		#1		read = 32'd3427522847;
		#1		read = 32'd3444701487;
		#1		read = 32'd3461750405;
		#1		read = 32'd3478667898;
		#1		read = 32'd3495452274;
		#1		read = 32'd3512101853;
		#1		read = 32'd3528614973;
		#1		read = 32'd3544989980;
		#1		read = 32'd3561225238;
		#1		read = 32'd3577319122;
		#1		read = 32'd3593270025;
		#1		read = 32'd3609076350;
		#1		read = 32'd3624736517;
		#1		read = 32'd3640248960;
		#1		read = 32'd3655612127;
		#1		read = 32'd3670824483;
		#1		read = 32'd3685884506;
		#1		read = 32'd3700790691;
		#1		read = 32'd3715541546;
		#1		read = 32'd3730135596;
		#1		read = 32'd3744571383;
		#1		read = 32'd3758847462;
		#1		read = 32'd3772962406;
		#1		read = 32'd3786914803;
		#1		read = 32'd3800703259;
		#1		read = 32'd3814326395;
		#1		read = 32'd3827782847;
		#1		read = 32'd3841071271;
		#1		read = 32'd3854190337;
		#1		read = 32'd3867138735;
		#1		read = 32'd3879915168;
		#1		read = 32'd3892518359;
		#1		read = 32'd3904947049;
		#1		read = 32'd3917199993;
		#1		read = 32'd3929275968;
		#1		read = 32'd3941173764;
		#1		read = 32'd3952892194;
		#1		read = 32'd3964430083;
		#1		read = 32'd3975786280;
		#1		read = 32'd3986959648;
		#1		read = 32'd3997949070;
		#1		read = 32'd4008753447;
		#1		read = 32'd4019371698;
		#1		read = 32'd4029802762;
		#1		read = 32'd4040045596;
		#1		read = 32'd4050099175;
		#1		read = 32'd4059962495;
		#1		read = 32'd4069634568;
		#1		read = 32'd4079114427;
		#1		read = 32'd4088401125;
		#1		read = 32'd4097493733;
		#1		read = 32'd4106391342;
		#1		read = 32'd4115093061;
		#1		read = 32'd4123598021;
		#1		read = 32'd4131905371;
		#1		read = 32'd4140014281;
		#1		read = 32'd4147923939;
		#1		read = 32'd4155633555;
		#1		read = 32'd4163142358;
		#1		read = 32'd4170449597;
		#1		read = 32'd4177554540;
		#1		read = 32'd4184456478;
		#1		read = 32'd4191154721;
		#1		read = 32'd4197648598;
		#1		read = 32'd4203937461;
		#1		read = 32'd4210020679;
		#1		read = 32'd4215897646;
		#1		read = 32'd4221567773;
		#1		read = 32'd4227030494;
		#1		read = 32'd4232285261;
		#1		read = 32'd4237331550;
		#1		read = 32'd4242168856;
		#1		read = 32'd4246796695;
		#1		read = 32'd4251214605;
		#1		read = 32'd4255422143;
		#1		read = 32'd4259418889;
		#1		read = 32'd4263204444;
		#1		read = 32'd4266778428;
		#1		read = 32'd4270140484;
		#1		read = 32'd4273290277;
		#1		read = 32'd4276227490;
		#1		read = 32'd4278951831;
		#1		read = 32'd4281463027;
		#1		read = 32'd4283760827;
		#1		read = 32'd4285845001;
		#1		read = 32'd4287715340;
		#1		read = 32'd4289371659;
		#1		read = 32'd4290813790;
		#1		read = 32'd4292041589;
		#1		read = 32'd4293054935;
		#1		read = 32'd4293853726;
		#1		read = 32'd4294437881;
		#1		read = 32'd4294807343;
		#1		read = 32'd4294962074;
		#1		read = 32'd4294902059;
		#1		read = 32'd4294627304;
		#1		read = 32'd4294137836;
		#1		read = 32'd4293433705;
		#1		read = 32'd4292514981;
		#1		read = 32'd4291381755;
		#1		read = 32'd4290034141;
		#1		read = 32'd4288472274;
		#1		read = 32'd4286696310;
		#1		read = 32'd4284706426;
		#1		read = 32'd4282502822;
		#1		read = 32'd4280085718;
		#1		read = 32'd4277455355;
		#1		read = 32'd4274611997;
		#1		read = 32'd4271555928;
		#1		read = 32'd4268287453;
		#1		read = 32'd4264806900;
		#1		read = 32'd4261114616;
		#1		read = 32'd4257210971;
		#1		read = 32'd4253096355;
		#1		read = 32'd4248771179;
		#1		read = 32'd4244235877;
		#1		read = 32'd4239490901;
		#1		read = 32'd4234536726;
		#1		read = 32'd4229373847;
		#1		read = 32'd4224002781;
		#1		read = 32'd4218424065;
		#1		read = 32'd4212638256;
		#1		read = 32'd4206645934;
		#1		read = 32'd4200447698;
		#1		read = 32'd4194044166;
		#1		read = 32'd4187435981;
		#1		read = 32'd4180623801;
		#1		read = 32'd4173608310;
		#1		read = 32'd4166390207;
		#1		read = 32'd4158970216;
		#1		read = 32'd4151349078;
		#1		read = 32'd4143527555;
		#1		read = 32'd4135506429;
		#1		read = 32'd4127286502;
		#1		read = 32'd4118868597;
		#1		read = 32'd4110253555;
		#1		read = 32'd4101442238;
		#1		read = 32'd4092435526;
		#1		read = 32'd4083234321;
		#1		read = 32'd4073839542;
		#1		read = 32'd4064252130;
		#1		read = 32'd4054473042;
		#1		read = 32'd4044503256;
		#1		read = 32'd4034343771;
		#1		read = 32'd4023995601;
		#1		read = 32'd4013459781;
		#1		read = 32'd4002737365;
		#1		read = 32'd3991829426;
		#1		read = 32'd3980737053;
		#1		read = 32'd3969461357;
		#1		read = 32'd3958003464;
		#1		read = 32'd3946364521;
		#1		read = 32'd3934545691;
		#1		read = 32'd3922548157;
		#1		read = 32'd3910373118;
		#1		read = 32'd3898021791;
		#1		read = 32'd3885495412;
		#1		read = 32'd3872795233;
		#1		read = 32'd3859922524;
		#1		read = 32'd3846878573;
		#1		read = 32'd3833664684;
		#1		read = 32'd3820282178;
		#1		read = 32'd3806732393;
		#1		read = 32'd3793016685;
		#1		read = 32'd3779136426;
		#1		read = 32'd3765093002;
		#1		read = 32'd3750887819;
		#1		read = 32'd3736522296;
		#1		read = 32'd3721997871;
		#1		read = 32'd3707315996;
		#1		read = 32'd3692478139;
		#1		read = 32'd3677485784;
		#1		read = 32'd3662340430;
		#1		read = 32'd3647043592;
		#1		read = 32'd3631596798;
		#1		read = 32'd3616001595;
		#1		read = 32'd3600259541;
		#1		read = 32'd3584372211;
		#1		read = 32'd3568341193;
		#1		read = 32'd3552168090;
		#1		read = 32'd3535854521;
		#1		read = 32'd3519402115;
		#1		read = 32'd3502812519;
		#1		read = 32'd3486087390;
		#1		read = 32'd3469228403;
		#1		read = 32'd3452237242;
		#1		read = 32'd3435115607;
		#1		read = 32'd3417865210;
		#1		read = 32'd3400487776;
		#1		read = 32'd3382985042;
		#1		read = 32'd3365358759;
		#1		read = 32'd3347610690;
		#1		read = 32'd3329742609;
		#1		read = 32'd3311756303;
		#1		read = 32'd3293653571;
		#1		read = 32'd3275436223;
		#1		read = 32'd3257106080;
		#1		read = 32'd3238664976;
		#1		read = 32'd3220114755;
		#1		read = 32'd3201457272;
		#1		read = 32'd3182694392;
		#1		read = 32'd3163827992;
		#1		read = 32'd3144859959;
		#1		read = 32'd3125792188;
		#1		read = 32'd3106626588;
		#1		read = 32'd3087365074;
		#1		read = 32'd3068009573;
		#1		read = 32'd3048562020;
		#1		read = 32'd3029024360;
		#1		read = 32'd3009398546;
		#1		read = 32'd2989686542;
		#1		read = 32'd2969890318;
		#1		read = 32'd2950011854;
		#1		read = 32'd2930053138;
		#1		read = 32'd2910016166;
		#1		read = 32'd2889902941;
		#1		read = 32'd2869715475;
		#1		read = 32'd2849455786;
		#1		read = 32'd2829125901;
		#1		read = 32'd2808727851;
		#1		read = 32'd2788263679;
		#1		read = 32'd2767735428;
		#1		read = 32'd2747145153;
		#1		read = 32'd2726494912;
		#1		read = 32'd2705786771;
		#1		read = 32'd2685022800;
		#1		read = 32'd2664205075;
		#1		read = 32'd2643335679;
		#1		read = 32'd2622416697;
		#1		read = 32'd2601450223;
		#1		read = 32'd2580438353;
		#1		read = 32'd2559383187;
		#1		read = 32'd2538286832;
		#1		read = 32'd2517151397;
		#1		read = 32'd2495978996;
		#1		read = 32'd2474771745;
		#1		read = 32'd2453531765;
		#1		read = 32'd2432261182;
		#1		read = 32'd2410962120;
		#1		read = 32'd2389636711;
		#1		read = 32'd2368287087;
		#1		read = 32'd2346915383;
		#1		read = 32'd2325523735;
		#1		read = 32'd2304114284;
		#1		read = 32'd2282689170;
		#1		read = 32'd2261250535;
		#1		read = 32'd2239800524;
		#1		read = 32'd2218341282;
		#1		read = 32'd2196874953;
		#1		read = 32'd2175403686;
		#1		read = 32'd2153929626;
		#1		read = 32'd2132454922;
		#1		read = 32'd2110981721;
		#1		read = 32'd2089512170;
		#1		read = 32'd2068048416;
		#1		read = 32'd2046592605;
		#1		read = 32'd2025146883;
		#1		read = 32'd2003713396;
		#1		read = 32'd1982294284;
		#1		read = 32'd1960891692;
		#1		read = 32'd1939507759;
		#1		read = 32'd1918144623;
		#1		read = 32'd1896804421;
		#1		read = 32'd1875489287;
		#1		read = 32'd1854201352;
		#1		read = 32'd1832942744;
		#1		read = 32'd1811715591;
		#1		read = 32'd1790522014;
		#1		read = 32'd1769364133;
		#1		read = 32'd1748244064;
		#1		read = 32'd1727163918;
		#1		read = 32'd1706125804;
		#1		read = 32'd1685131826;
		#1		read = 32'd1664184082;
		#1		read = 32'd1643284667;
		#1		read = 32'd1622435673;
		#1		read = 32'd1601639182;
		#1		read = 32'd1580897276;
		#1		read = 32'd1560212027;
		#1		read = 32'd1539585506;
		#1		read = 32'd1519019773;
		#1		read = 32'd1498516887;
		#1		read = 32'd1478078897;
		#1		read = 32'd1457707846;
		#1		read = 32'd1437405773;
		#1		read = 32'd1417174707;
		#1		read = 32'd1397016671;
		#1		read = 32'd1376933681;
		#1		read = 32'd1356927745;
		#1		read = 32'd1337000865;
		#1		read = 32'd1317155032;
		#1		read = 32'd1297392231;
		#1		read = 32'd1277714439;
		#1		read = 32'd1258123623;
		#1		read = 32'd1238621742;
		#1		read = 32'd1219210746;
		#1		read = 32'd1199892577;
		#1		read = 32'd1180669167;
		#1		read = 32'd1161542437;
		#1		read = 32'd1142514300;
		#1		read = 32'd1123586659;
		#1		read = 32'd1104761408;
		#1		read = 32'd1086040427;
		#1		read = 32'd1067425590;
		#1		read = 32'd1048918758;
		#1		read = 32'd1030521782;
		#1		read = 32'd1012236501;
		#1		read = 32'd994064743;
		#1		read = 32'd976008327;
		#1		read = 32'd958069057;
		#1		read = 32'd940248727;
		#1		read = 32'd922549120;
		#1		read = 32'd904972006;
		#1		read = 32'd887519141;
		#1		read = 32'd870192272;
		#1		read = 32'd852993131;
		#1		read = 32'd835923438;
		#1		read = 32'd818984900;
		#1		read = 32'd802179211;
		#1		read = 32'd785508051;
		#1		read = 32'd768973087;
		#1		read = 32'd752575974;
		#1		read = 32'd736318349;
		#1		read = 32'd720201841;
		#1		read = 32'd704228059;
		#1		read = 32'd688398602;
		#1		read = 32'd672715052;
		#1		read = 32'd657178977;
		#1		read = 32'd641791932;
		#1		read = 32'd626555455;
		#1		read = 32'd611471069;
		#1		read = 32'd596540283;
		#1		read = 32'd581764591;
		#1		read = 32'd567145468;
		#1		read = 32'd552684379;
		#1		read = 32'd538382768;
		#1		read = 32'd524242066;
		#1		read = 32'd510263686;
		#1		read = 32'd496449027;
		#1		read = 32'd482799471;
		#1		read = 32'd469316381;
		#1		read = 32'd456001106;
		#1		read = 32'd442854979;
		#1		read = 32'd429879313;
		#1		read = 32'd417075406;
		#1		read = 32'd404444538;
		#1		read = 32'd391987973;
		#1		read = 32'd379706956;
		#1		read = 32'd367602715;
		#1		read = 32'd355676460;
		#1		read = 32'd343929385;
		#1		read = 32'd332362664;
		#1		read = 32'd320977453;
		#1		read = 32'd309774892;
		#1		read = 32'd298756100;
		#1		read = 32'd287922179;
		#1		read = 32'd277274213;
		#1		read = 32'd266813266;
		#1		read = 32'd256540384;
		#1		read = 32'd246456595;
		#1		read = 32'd236562908;
		#1		read = 32'd226860311;
		#1		read = 32'd217349774;
		#1		read = 32'd208032250;
		#1		read = 32'd198908668;
		#1		read = 32'd189979943;
		#1		read = 32'd181246967;
		#1		read = 32'd172710612;
		#1		read = 32'd164371733;
		#1		read = 32'd156231164;
		#1		read = 32'd148289719;
		#1		read = 32'd140548191;
		#1		read = 32'd133007354;
		#1		read = 32'd125667964;
		#1		read = 32'd118530754;
		#1		read = 32'd111596437;
		#1		read = 32'd104865708;
		#1		read = 32'd98339238;
		#1		read = 32'd92017682;
		#1		read = 32'd85901670;
		#1		read = 32'd79991814;
		#1		read = 32'd74288706;
		#1		read = 32'd68792916;
		#1		read = 32'd63504993;
		#1		read = 32'd58425466;
		#1		read = 32'd53554844;
		#1		read = 32'd48893612;
		#1		read = 32'd44442238;
		#1		read = 32'd40201166;
		#1		read = 32'd36170821;
		#1		read = 32'd32351605;
		#1		read = 32'd28743900;
		#1		read = 32'd25348068;
		#1		read = 32'd22164448;
		#1		read = 32'd19193358;
		#1		read = 32'd16435095;
		#1		read = 32'd13889935;
		#1		read = 32'd11558132;
		#1		read = 32'd9439921;
		#1		read = 32'd7535512;
		#1		read = 32'd5845096;
		#1		read = 32'd4368842;
		#1		read = 32'd3106898;
		#1		read = 32'd2059389;
		#1		read = 32'd1226422;
		#1		read = 32'd608078;
		#1		read = 32'd204420;
		#1		read = 32'd15488;
		#1		read = 32'd41301;
		#1		read = 32'd281857;
		#1		read = 32'd737131;
		#1		read = 32'd1407078;
		#1		read = 32'd2291631;
		#1		read = 32'd3390701;
		#1		read = 32'd4704179;
		#1		read = 32'd6231933;
		#1		read = 32'd7973810;
		#1		read = 32'd9929636;
		#1		read = 32'd12099216;
		#1		read = 32'd14482333;
		#1		read = 32'd17078748;
		#1		read = 32'd19888202;
		#1		read = 32'd22910413;
		#1		read = 32'd26145081;
		#1		read = 32'd29591880;
		#1		read = 32'd33250466;
		#1		read = 32'd37120475;
		#1		read = 32'd41201517;
		#1		read = 32'd45493187;
		#1		read = 32'd49995053;
		#1		read = 32'd54706667;
		#1		read = 32'd59627556;
		#1		read = 32'd64757230;
		#1		read = 32'd70095174;
		#1		read = 32'd75640855;
		#1		read = 32'd81393719;
		#1		read = 32'd87353191;
		#1		read = 32'd93518673;
		#1		read = 32'd99889551;
		#1		read = 32'd106465186;
		#1		read = 32'd113244921;
		#1		read = 32'd120228078;
		#1		read = 32'd127413960;
		#1		read = 32'd134801846;
		#1		read = 32'd142390999;
		#1		read = 32'd150180660;
		#1		read = 32'd158170049;
		#1		read = 32'd166358368;
		#1		read = 32'd174744798;
		#1		read = 32'd183328500;
		#1		read = 32'd192108616;
		#1		read = 32'd201084268;
		#1		read = 32'd210254558;
		#1		read = 32'd219618570;
		#1		read = 32'd229175366;
		#1		read = 32'd238923992;
		#1		read = 32'd248863472;
		#1		read = 32'd258992812;
		#1		read = 32'd269311000;
		#1		read = 32'd279817004;
		#1		read = 32'd290509772;
		#1		read = 32'd301388237;
		#1		read = 32'd312451310;
		#1		read = 32'd323697884;
		#1		read = 32'd335126835;
		#1		read = 32'd346737021;
		#1		read = 32'd358527279;
		#1		read = 32'd370496432;
		#1		read = 32'd382643282;
		#1		read = 32'd394966615;
		#1		read = 32'd407465198;
		#1		read = 32'd420137781;
		#1		read = 32'd432983097;
		#1		read = 32'd445999862;
		#1		read = 32'd459186774;
		#1		read = 32'd472542515;
		#1		read = 32'd486065748;
		#1		read = 32'd499755121;
		#1		read = 32'd513609266;
		#1		read = 32'd527626797;
		#1		read = 32'd541806312;
		#1		read = 32'd556146394;
		#1		read = 32'd570645608;
		#1		read = 32'd585302505;
		#1		read = 32'd600115618;
		#1		read = 32'd615083467;
		#1		read = 32'd630204554;
		#1		read = 32'd645477369;
		#1		read = 32'd660900382;
		#1		read = 32'd676472053;
		#1		read = 32'd692190824;
		#1		read = 32'd708055123;
		#1		read = 32'd724063363;
		#1		read = 32'd740213944;
		#1		read = 32'd756505251;
		#1		read = 32'd772935655;
		#1		read = 32'd789503512;
		#1		read = 32'd806207167;
		#1		read = 32'd823044948;
		#1		read = 32'd840015171;
		#1		read = 32'd857116140;
		#1		read = 32'd874346145;
		#1		read = 32'd891703463;
		#1		read = 32'd909186358;
		#1		read = 32'd926793081;
		#1		read = 32'd944521873;
		#1		read = 32'd962370959;
		#1		read = 32'd980338556;
		#1		read = 32'd998422866;
		#1		read = 32'd1016622082;
		#1		read = 32'd1034934383;
		#1		read = 32'd1053357937;
		#1		read = 32'd1071890904;
		#1		read = 32'd1090531428;
		#1		read = 32'd1109277647;
		#1		read = 32'd1128127686;
		#1		read = 32'd1147079660;
		#1		read = 32'd1166131673;
		#1		read = 32'd1185281821;
		#1		read = 32'd1204528187;
		#1		read = 32'd1223868849;
		#1		read = 32'd1243301872;
		#1		read = 32'd1262825311;
		#1		read = 32'd1282437216;
		#1		read = 32'd1302135625;
		#1		read = 32'd1321918568;
		#1		read = 32'd1341784067;
		#1		read = 32'd1361730135;
		#1		read = 32'd1381754777;
		#1		read = 32'd1401855992;
		#1		read = 32'd1422031770;
		#1		read = 32'd1442280091;
		#1		read = 32'd1462598933;
		#1		read = 32'd1482986262;
		#1		read = 32'd1503440041;
		#1		read = 32'd1523958223;
		#1		read = 32'd1544538757;
		#1		read = 32'd1565179586;
		#1		read = 32'd1585878644;
		#1		read = 32'd1606633862;
		#1		read = 32'd1627443165;
		#1		read = 32'd1648304472;
		#1		read = 32'd1669215696;
		#1		read = 32'd1690174746;
		#1		read = 32'd1711179527;
		#1		read = 32'd1732227938;
		#1		read = 32'd1753317874;
		#1		read = 32'd1774447227;
		#1		read = 32'd1795613882;
		#1		read = 32'd1816815725;
		#1		read = 32'd1838050634;
		#1		read = 32'd1859316486;
		#1		read = 32'd1880611154;
		#1		read = 32'd1901932510;
		#1		read = 32'd1923278420;
		#1		read = 32'd1944646751;
		#1		read = 32'd1966035365;
		#1		read = 32'd1987442124;
		#1		read = 32'd2008864887;
		#1		read = 32'd2030301512;
		#1		read = 32'd2051749854;
		#1		read = 32'd2073207771;
		#1		read = 32'd2094673114;
		#1		read = 32'd2116143739;
		#1		read = 32'd2137617497;
		#1		read = 32'd2159092243;
		#1		read = 32'd2180565827;
		#1		read = 32'd2202036103;
		#1		read = 32'd2223500924;
		#1		read = 32'd2244958144;
		#1		read = 32'd2266405616;
		#1		read = 32'd2287841195;
		#1		read = 32'd2309262740;
		#1		read = 32'd2330668106;
		#1		read = 32'd2352055154;
		#1		read = 32'd2373421745;
		#1		read = 32'd2394765743;
		#1		read = 32'd2416085013;
		#1		read = 32'd2437377422;
		#1		read = 32'd2458640843;
		#1		read = 32'd2479873148;
		#1		read = 32'd2501072214;
		#1		read = 32'd2522235922;
		#1		read = 32'd2543362155;
		#1		read = 32'd2564448800;
		#1		read = 32'd2585493749;
		#1		read = 32'd2606494898;
		#1		read = 32'd2627450146;
		#1		read = 32'd2648357397;
		#1		read = 32'd2669214562;
		#1		read = 32'd2690019554;
		#1		read = 32'd2710770293;
		#1		read = 32'd2731464703;
		#1		read = 32'd2752100716;
		#1		read = 32'd2772676268;
		#1		read = 32'd2793189301;
		#1		read = 32'd2813637764;
		#1		read = 32'd2834019612;
		#1		read = 32'd2854332808;
		#1		read = 32'd2874575318;
		#1		read = 32'd2894745121;
		#1		read = 32'd2914840197;
		#1		read = 32'd2934858539;
		#1		read = 32'd2954798144;
		#1		read = 32'd2974657018;
		#1		read = 32'd2994433176;
		#1		read = 32'd3014124639;
		#1		read = 32'd3033729439;
		#1		read = 32'd3053245615;
		#1		read = 32'd3072671215;
		#1		read = 32'd3092004298;
		#1		read = 32'd3111242929;
		#1		read = 32'd3130385185;
		#1		read = 32'd3149429152;
		#1		read = 32'd3168372925;
		#1		read = 32'd3187214610;
		#1		read = 32'd3205952323;
		#1		read = 32'd3224584190;
		#1		read = 32'd3243108348;
		#1		read = 32'd3261522944;
		#1		read = 32'd3279826137;
		#1		read = 32'd3298016097;
		#1		read = 32'd3316091004;
		#1		read = 32'd3334049052;
		#1		read = 32'd3351888444;
		#1		read = 32'd3369607397;
		#1		read = 32'd3387204138;
		#1		read = 32'd3404676909;
		#1		read = 32'd3422023961;
		#1		read = 32'd3439243560;
		#1		read = 32'd3456333984;
		#1		read = 32'd3473293524;
		#1		read = 32'd3490120485;
		#1		read = 32'd3506813182;
		#1		read = 32'd3523369948;
		#1		read = 32'd3539789127;
		#1		read = 32'd3556069076;
		#1		read = 32'd3572208168;
		#1		read = 32'd3588204788;
		#1		read = 32'd3604057338;
		#1		read = 32'd3619764231;
		#1		read = 32'd3635323898;
		#1		read = 32'd3650734782;
		#1		read = 32'd3665995341;
		#1		read = 32'd3681104052;
		#1		read = 32'd3696059401;
		#1		read = 32'd3710859894;
		#1		read = 32'd3725504050;
		#1		read = 32'd3739990406;
		#1		read = 32'd3754317513;
		#1		read = 32'd3768483938;
		#1		read = 32'd3782488263;
		#1		read = 32'd3796329090;
		#1		read = 32'd3810005034;
		#1		read = 32'd3823514727;
		#1		read = 32'd3836856818;
		#1		read = 32'd3850029973;
		#1		read = 32'd3863032875;
		#1		read = 32'd3875864223;
		#1		read = 32'd3888522735;
		#1		read = 32'd3901007145;
		#1		read = 32'd3913316203;
		#1		read = 32'd3925448680;
		#1		read = 32'd3937403362;
		#1		read = 32'd3949179053;
		#1		read = 32'd3960774576;
		#1		read = 32'd3972188772;
		#1		read = 32'd3983420499;
		#1		read = 32'd3994468633;
		#1		read = 32'd4005332071;
		#1		read = 32'd4016009725;
		#1		read = 32'd4026500528;
		#1		read = 32'd4036803431;
		#1		read = 32'd4046917404;
		#1		read = 32'd4056841435;
		#1		read = 32'd4066574531;
		#1		read = 32'd4076115721;
		#1		read = 32'd4085464048;
		#1		read = 32'd4094618579;
		#1		read = 32'd4103578399;
		#1		read = 32'd4112342610;
		#1		read = 32'd4120910337;
		#1		read = 32'd4129280723;
		#1		read = 32'd4137452932;
		#1		read = 32'd4145426144;
		#1		read = 32'd4153199565;
		#1		read = 32'd4160772415;
		#1		read = 32'd4168143938;
		#1		read = 32'd4175313397;
		#1		read = 32'd4182280075;
		#1		read = 32'd4189043274;
		#1		read = 32'd4195602319;
		#1		read = 32'd4201956555;
		#1		read = 32'd4208105344;
		#1		read = 32'd4214048073;
		#1		read = 32'd4219784148;
		#1		read = 32'd4225312994;
		#1		read = 32'd4230634059;
		#1		read = 32'd4235746810;
		#1		read = 32'd4240650737;
		#1		read = 32'd4245345349;
		#1		read = 32'd4249830177;
		#1		read = 32'd4254104771;
		#1		read = 32'd4258168706;
		#1		read = 32'd4262021573;
		#1		read = 32'd4265662989;
		#1		read = 32'd4269092588;
		#1		read = 32'd4272310029;
		#1		read = 32'd4275314988;
		#1		read = 32'd4278107166;
		#1		read = 32'd4280686283;
		#1		read = 32'd4283052082;
		#1		read = 32'd4285204326;
		#1		read = 32'd4287142800;
		#1		read = 32'd4288867310;
		#1		read = 32'd4290377682;
		#1		read = 32'd4291673768;
		#1		read = 32'd4292755436;
		#1		read = 32'd4293622578;
		#1		read = 32'd4294275109;
		#1		read = 32'd4294712962;
		#1		read = 32'd4294936094;
		#1		read = 32'd4294944483;
		#1		read = 32'd4294738127;
		#1		read = 32'd4294317048;
		#1		read = 32'd4293681287;
		#1		read = 32'd4292830908;
		#1		read = 32'd4291765996;
		#1		read = 32'd4290486658;
		#1		read = 32'd4288993021;
		#1		read = 32'd4287285236;
		#1		read = 32'd4285363471;
		#1		read = 32'd4283227921;
		#1		read = 32'd4280878798;
		#1		read = 32'd4278316337;
		#1		read = 32'd4275540794;
		#1		read = 32'd4272552448;
		#1		read = 32'd4269351597;
		#1		read = 32'd4265938560;
		#1		read = 32'd4262313680;
		#1		read = 32'd4258477319;
		#1		read = 32'd4254429860;
		#1		read = 32'd4250171708;
		#1		read = 32'd4245703289;
		#1		read = 32'd4241025050;
		#1		read = 32'd4236137458;
		#1		read = 32'd4231041003;
		#1		read = 32'd4225736194;
		#1		read = 32'd4220223561;
		#1		read = 32'd4214503656;
		#1		read = 32'd4208577051;
		#1		read = 32'd4202444338;
		#1		read = 32'd4196106131;
		#1		read = 32'd4189563063;
		#1		read = 32'd4182815789;
		#1		read = 32'd4175864983;
		#1		read = 32'd4168711341;
		#1		read = 32'd4161355578;
		#1		read = 32'd4153798430;
		#1		read = 32'd4146040651;
		#1		read = 32'd4138083019;
		#1		read = 32'd4129926328;
		#1		read = 32'd4121571395;
		#1		read = 32'd4113019055;
		#1		read = 32'd4104270162;
		#1		read = 32'd4095325593;
		#1		read = 32'd4086186241;
		#1		read = 32'd4076853020;
		#1		read = 32'd4067326864;
		#1		read = 32'd4057608726;
		#1		read = 32'd4047699576;
		#1		read = 32'd4037600407;
		#1		read = 32'd4027312227;
		#1		read = 32'd4016836066;
		#1		read = 32'd4006172971;
		#1		read = 32'd3995324009;
		#1		read = 32'd3984290265;
		#1		read = 32'd3973072841;
		#1		read = 32'd3961672860;
		#1		read = 32'd3950091462;
		#1		read = 32'd3938329804;
		#1		read = 32'd3926389063;
		#1		read = 32'd3914270433;
		#1		read = 32'd3901975126;
		#1		read = 32'd3889504371;
		#1		read = 32'd3876859416;
		#1		read = 32'd3864041524;
		#1		read = 32'd3851051979;
		#1		read = 32'd3837892077;
		#1		read = 32'd3824563136;
		#1		read = 32'd3811066489;
		#1		read = 32'd3797403485;
		#1		read = 32'd3783575490;
		#1		read = 32'd3769583887;
		#1		read = 32'd3755430076;
		#1		read = 32'd3741115472;
		#1		read = 32'd3726641505;
		#1		read = 32'd3712009624;
		#1		read = 32'd3697221292;
		#1		read = 32'd3682277987;
		#1		read = 32'd3667181204;
		#1		read = 32'd3651932453;
		#1		read = 32'd3636533258;
		#1		read = 32'd3620985159;
		#1		read = 32'd3605289712;
		#1		read = 32'd3589448485;
		#1		read = 32'd3573463062;
		#1		read = 32'd3557335043;
		#1		read = 32'd3541066040;
		#1		read = 32'd3524657680;
		#1		read = 32'd3508111604;
		#1		read = 32'd3491429466;
		#1		read = 32'd3474612934;
		#1		read = 32'd3457663691;
		#1		read = 32'd3440583431;
		#1		read = 32'd3423373862;
		#1		read = 32'd3406036705;
		#1		read = 32'd3388573693;
		#1		read = 32'd3370986574;
		#1		read = 32'd3353277106;
		#1		read = 32'd3335447059;
		#1		read = 32'd3317498216;
		#1		read = 32'd3299432374;
		#1		read = 32'd3281251337;
		#1		read = 32'd3262956925;
		#1		read = 32'd3244550966;
		#1		read = 32'd3226035301;
		#1		read = 32'd3207411782;
		#1		read = 32'd3188682271;
		#1		read = 32'd3169848641;
		#1		read = 32'd3150912776;
		#1		read = 32'd3131876568;
		#1		read = 32'd3112741922;
		#1		read = 32'd3093510751;
		#1		read = 32'd3074184978;
		#1		read = 32'd3054766536;
		#1		read = 32'd3035257366;
		#1		read = 32'd3015659419;
		#1		read = 32'd2995974656;
		#1		read = 32'd2976205044;
		#1		read = 32'd2956352561;
		#1		read = 32'd2936419191;
		#1		read = 32'd2916406929;
		#1		read = 32'd2896317775;
		#1		read = 32'd2876153738;
		#1		read = 32'd2855916835;
		#1		read = 32'd2835609089;
		#1		read = 32'd2815232531;
		#1		read = 32'd2794789199;
		#1		read = 32'd2774281136;
		#1		read = 32'd2753710395;
		#1		read = 32'd2733079031;
		#1		read = 32'd2712389108;
		#1		read = 32'd2691642696;
		#1		read = 32'd2670841867;
		#1		read = 32'd2649988704;
		#1		read = 32'd2629085290;
		#1		read = 32'd2608133716;
		#1		read = 32'd2587136078;
		#1		read = 32'd2566094475;
		#1		read = 32'd2545011012;
		#1		read = 32'd2523887796;
		#1		read = 32'd2502726939;
		#1		read = 32'd2481530559;
		#1		read = 32'd2460300774;
		#1		read = 32'd2439039708;
		#1		read = 32'd2417749487;
		#1		read = 32'd2396432239;
		#1		read = 32'd2375090096;
		#1		read = 32'd2353725193;
		#1		read = 32'd2332339666;
		#1		read = 32'd2310935654;
		#1		read = 32'd2289515297;
		#1		read = 32'd2268080736;
		#1		read = 32'd2246634116;
		#1		read = 32'd2225177581;
		#1		read = 32'd2203713277;
		#1		read = 32'd2182243349;
		#1		read = 32'd2160769946;
		#1		read = 32'd2139295214;
		#1		read = 32'd2117821301;
		#1		read = 32'd2096350354;
		#1		read = 32'd2074884521;
		#1		read = 32'd2053425947;
		#1		read = 32'd2031976779;
		#1		read = 32'd2010539162;
		#1		read = 32'd1989115239;
		#1		read = 32'd1967707152;
		#1		read = 32'd1946317043;
		#1		read = 32'd1924947051;
		#1		read = 32'd1903599312;
		#1		read = 32'd1882275961;
		#1		read = 32'd1860979131;
		#1		read = 32'd1839710951;
		#1		read = 32'd1818473548;
		#1		read = 32'd1797269046;
		#1		read = 32'd1776099565;
		#1		read = 32'd1754967222;
		#1		read = 32'd1733874131;
		#1		read = 32'd1712822400;
		#1		read = 32'd1691814135;
		#1		read = 32'd1670851436;
		#1		read = 32'd1649936400;
		#1		read = 32'd1629071119;
		#1		read = 32'd1608257678;
		#1		read = 32'd1587498160;
		#1		read = 32'd1566794639;
		#1		read = 32'd1546149187;
		#1		read = 32'd1525563868;
		#1		read = 32'd1505040740;
		#1		read = 32'd1484581857;
		#1		read = 32'd1464189262;
		#1		read = 32'd1443864997;
		#1		read = 32'd1423611093;
		#1		read = 32'd1403429575;
		#1		read = 32'd1383322463;
		#1		read = 32'd1363291766;
		#1		read = 32'd1343339487;
		#1		read = 32'd1323467622;
		#1		read = 32'd1303678158;
		#1		read = 32'd1283973074;
		#1		read = 32'd1264354340;
		#1		read = 32'd1244823918;
		#1		read = 32'd1225383762;
		#1		read = 32'd1206035815;
		#1		read = 32'd1186782012;
		#1		read = 32'd1167624278;
		#1		read = 32'd1148564529;
		#1		read = 32'd1129604672;
		#1		read = 32'd1110746601;
		#1		read = 32'd1091992203;
		#1		read = 32'd1073343354;
		#1		read = 32'd1054801918;
		#1		read = 32'd1036369749;
		#1		read = 32'd1018048690;
		#1		read = 32'd999840574;
		#1		read = 32'd981747221;
		#1		read = 32'd963770441;
		#1		read = 32'd945912032;
		#1		read = 32'd928173778;
		#1		read = 32'd910557455;
		#1		read = 32'd893064823;
		#1		read = 32'd875697632;
		#1		read = 32'd858457618;
		#1		read = 32'd841346506;
		#1		read = 32'd824366007;
		#1		read = 32'd807517818;
		#1		read = 32'd790803625;
		#1		read = 32'd774225098;
		#1		read = 32'd757783896;
		#1		read = 32'd741481664;
		#1		read = 32'd725320030;
		#1		read = 32'd709300611;
		#1		read = 32'd693425009;
		#1		read = 32'd677694812;
		#1		read = 32'd662111593;
		#1		read = 32'd646676910;
		#1		read = 32'd631392306;
		#1		read = 32'd616259310;
		#1		read = 32'd601279435;
		#1		read = 32'd586454179;
		#1		read = 32'd571785025;
		#1		read = 32'd557273440;
		#1		read = 32'd542920874;
		#1		read = 32'd528728763;
		#1		read = 32'd514698526;
		#1		read = 32'd500831567;
		#1		read = 32'd487129271;
		#1		read = 32'd473593009;
		#1		read = 32'd460224135;
		#1		read = 32'd447023986;
		#1		read = 32'd433993881;
		#1		read = 32'd421135123;
		#1		read = 32'd408448999;
		#1		read = 32'd395936778;
		#1		read = 32'd383599709;
		#1		read = 32'd371439027;
		#1		read = 32'd359455948;
		#1		read = 32'd347651671;
		#1		read = 32'd336027375;
		#1		read = 32'd324584223;
		#1		read = 32'd313323360;
		#1		read = 32'd302245911;
		#1		read = 32'd291352984;
		#1		read = 32'd280645669;
		#1		read = 32'd270125036;
		#1		read = 32'd259792138;
		#1		read = 32'd249648007;
		#1		read = 32'd239693658;
		#1		read = 32'd229930086;
		#1		read = 32'd220358269;
		#1		read = 32'd210979162;
		#1		read = 32'd201793704;
		#1		read = 32'd192802813;
		#1		read = 32'd184007389;
		#1		read = 32'd175408311;
		#1		read = 32'd167006438;
		#1		read = 32'd158802612;
		#1		read = 32'd150797652;
		#1		read = 32'd142992360;
		#1		read = 32'd135387514;
		#1		read = 32'd127983877;
		#1		read = 32'd120782188;
		#1		read = 32'd113783167;
		#1		read = 32'd106987514;
		#1		read = 32'd100395910;
		#1		read = 32'd94009013;
		#1		read = 32'd87827461;
		#1		read = 32'd81851873;
		#1		read = 32'd76082847;
		#1		read = 32'd70520959;
		#1		read = 32'd65166766;
		#1		read = 32'd60020802;
		#1		read = 32'd55083583;
		#1		read = 32'd50355603;
		#1		read = 32'd45837333;
		#1		read = 32'd41529227;
		#1		read = 32'd37431714;
		#1		read = 32'd33545204;
		#1		read = 32'd29870087;
		#1		read = 32'd26406729;
		#1		read = 32'd23155477;
		#1		read = 32'd20116656;
		#1		read = 32'd17290570;
		#1		read = 32'd14677501;
		#1		read = 32'd12277712;
		#1		read = 32'd10091441;
		#1		read = 32'd8118908;
		#1		read = 32'd6360309;
		#1		read = 32'd4815821;
		#1		read = 32'd3485598;
		#1		read = 32'd2369773;
		#1		read = 32'd1468457;
		#1		read = 32'd781741;
		#1		read = 32'd309694;
		#1		read = 32'd52362;
		#1		read = 32'd9772;
		#1		read = 32'd181927;
		#1		read = 32'd568810;
		#1		read = 32'd1170384;
		#1		read = 32'd1986586;
		#1		read = 32'd3017337;
		#1		read = 32'd4262533;
		#1		read = 32'd5722049;
		#1		read = 32'd7395739;
		#1		read = 32'd9283436;
		#1		read = 32'd11384952;
		#1		read = 32'd13700075;
		#1		read = 32'd16228575;
		#1		read = 32'd18970199;
		#1		read = 32'd21924673;
		#1		read = 32'd25091700;
		#1		read = 32'd28470965;
		#1		read = 32'd32062130;
		#1		read = 32'd35864835;
		#1		read = 32'd39878700;
		#1		read = 32'd44103324;
		#1		read = 32'd48538284;
		#1		read = 32'd53183136;
		#1		read = 32'd58037418;
		#1		read = 32'd63100642;
		#1		read = 32'd68372302;
		#1		read = 32'd73851872;
		#1		read = 32'd79538804;
		#1		read = 32'd85432528;
		#1		read = 32'd91532455;
		#1		read = 32'd97837976;
		#1		read = 32'd104348460;
		#1		read = 32'd111063256;
		#1		read = 32'd117981692;
		#1		read = 32'd125103076;
		#1		read = 32'd132426697;
		#1		read = 32'd139951822;
		#1		read = 32'd147677699;
		#1		read = 32'd155603554;
		#1		read = 32'd163728596;
		#1		read = 32'd172052011;
		#1		read = 32'd180572968;
		#1		read = 32'd189290615;
		#1		read = 32'd198204079;
		#1		read = 32'd207312470;
		#1		read = 32'd216614876;
		#1		read = 32'd226110367;
		#1		read = 32'd235797994;
		#1		read = 32'd245676788;
		#1		read = 32'd255745761;
		#1		read = 32'd266003906;
		#1		read = 32'd276450198;
		#1		read = 32'd287083591;
		#1		read = 32'd297903023;
		#1		read = 32'd308907412;
		#1		read = 32'd320095656;
		#1		read = 32'd331466638;
		#1		read = 32'd343019220;
		#1		read = 32'd354752247;
		#1		read = 32'd366664546;
		#1		read = 32'd378754925;
		#1		read = 32'd391022175;
		#1		read = 32'd403465070;
		#1		read = 32'd416082366;
		#1		read = 32'd428872800;
		#1		read = 32'd441835094;
		#1		read = 32'd454967951;
		#1		read = 32'd468270058;
		#1		read = 32'd481740086;
		#1		read = 32'd495376686;
		#1		read = 32'd509178496;
		#1		read = 32'd523144135;
		#1		read = 32'd537272206;
		#1		read = 32'd551561297;
		#1		read = 32'd566009979;
		#1		read = 32'd580616808;
		#1		read = 32'd595380321;
		#1		read = 32'd610299044;
		#1		read = 32'd625371484;
		#1		read = 32'd640596133;
		#1		read = 32'd655971471;
		#1		read = 32'd671495958;
		#1		read = 32'd687168042;
		#1		read = 32'd702986158;
		#1		read = 32'd718948721;
		#1		read = 32'd735054137;
		#1		read = 32'd751300795;
		#1		read = 32'd767687070;
		#1		read = 32'd784211323;
		#1		read = 32'd800871902;
		#1		read = 32'd817667142;
		#1		read = 32'd834595362;
		#1		read = 32'd851654870;
		#1		read = 32'd868843959;
		#1		read = 32'd886160912;
		#1		read = 32'd903603995;
		#1		read = 32'd921171466;
		#1		read = 32'd938861567;
		#1		read = 32'd956672529;
		#1		read = 32'd974602571;
		#1		read = 32'd992649900;
		#1		read = 32'd1010812712;
		#1		read = 32'd1029089190;
		#1		read = 32'd1047477506;
		#1		read = 32'd1065975822;
		#1		read = 32'd1084582288;
		#1		read = 32'd1103295043;
		#1		read = 32'd1122112216;
		#1		read = 32'd1141031926;
		#1		read = 32'd1160052280;
		#1		read = 32'd1179171376;
		#1		read = 32'd1198387302;
		#1		read = 32'd1217698138;
		#1		read = 32'd1237101951;
		#1		read = 32'd1256596801;
		#1		read = 32'd1276180740;
		#1		read = 32'd1295851808;
		#1		read = 32'd1315608038;
		#1		read = 32'd1335447456;
		#1		read = 32'd1355368076;
		#1		read = 32'd1375367907;
		#1		read = 32'd1395444949;
		#1		read = 32'd1415597195;
		#1		read = 32'd1435822628;
		#1		read = 32'd1456119227;
		#1		read = 32'd1476484962;
		#1		read = 32'd1496917796;
		#1		read = 32'd1517415686;
		#1		read = 32'd1537976583;
		#1		read = 32'd1558598429;
		#1		read = 32'd1579279164;
		#1		read = 32'd1600016719;
		#1		read = 32'd1620809020;
		#1		read = 32'd1641653987;
		#1		read = 32'd1662549538;
		#1		read = 32'd1683493581;
		#1		read = 32'd1704484023;
		#1		read = 32'd1725518765;
		#1		read = 32'd1746595703;
		#1		read = 32'd1767712729;
		#1		read = 32'd1788867732;
		#1		read = 32'd1810058597;
		#1		read = 32'd1831283203;
		#1		read = 32'd1852539429;
		#1		read = 32'd1873825150;
		#1		read = 32'd1895138236;
		#1		read = 32'd1916476557;
		#1		read = 32'd1937837978;
		#1		read = 32'd1959220363;
		#1		read = 32'd1980621574;
		#1		read = 32'd2002039472;
		#1		read = 32'd2023471914;
		#1		read = 32'd2044916757;
		#1		read = 32'd2066371857;
		#1		read = 32'd2087835067;
		#1		read = 32'd2109304243;
		#1		read = 32'd2130777236;
		#1		read = 32'd2152251900;
		#1		read = 32'd2173726087;
		#1		read = 32'd2195197650;
		#1		read = 32'd2216664442;
		#1		read = 32'd2238124316;
		#1		read = 32'd2259575125;
		#1		read = 32'd2281014726;
		#1		read = 32'd2302440973;
		#1		read = 32'd2323851725;
		#1		read = 32'd2345244841;
		#1		read = 32'd2366618180;
		#1		read = 32'd2387969606;
		#1		read = 32'd2409296984;
		#1		read = 32'd2430598180;
		#1		read = 32'd2451871066;
		#1		read = 32'd2473113513;
		#1		read = 32'd2494323397;
		#1		read = 32'd2515498597;
		#1		read = 32'd2536636997;
		#1		read = 32'd2557736481;
		#1		read = 32'd2578794940;
		#1		read = 32'd2599810269;
		#1		read = 32'd2620780365;
		#1		read = 32'd2641703132;
		#1		read = 32'd2662576477;
		#1		read = 32'd2683398314;
		#1		read = 32'd2704166560;
		#1		read = 32'd2724879137;
		#1		read = 32'd2745533976;
		#1		read = 32'd2766129010;
		#1		read = 32'd2786662180;
		#1		read = 32'd2807131433;
		#1		read = 32'd2827534722;
		#1		read = 32'd2847870006;
		#1		read = 32'd2868135252;
		#1		read = 32'd2888328433;
		#1		read = 32'd2908447531;
		#1		read = 32'd2928490533;
		#1		read = 32'd2948455434;
		#1		read = 32'd2968340240;
		#1		read = 32'd2988142960;
		#1		read = 32'd3007861615;
		#1		read = 32'd3027494233;
		#1		read = 32'd3047038851;
		#1		read = 32'd3066493514;
		#1		read = 32'd3085856276;
		#1		read = 32'd3105125202;
		#1		read = 32'd3124298365;
		#1		read = 32'd3143373847;
		#1		read = 32'd3162349741;
		#1		read = 32'd3181224150;
		#1		read = 32'd3199995185;
		#1		read = 32'd3218660969;
		#1		read = 32'd3237219637;
		#1		read = 32'd3255669333;
		#1		read = 32'd3274008210;
		#1		read = 32'd3292234436;
		#1		read = 32'd3310346188;
		#1		read = 32'd3328341655;
		#1		read = 32'd3346219037;
		#1		read = 32'd3363976546;
		#1		read = 32'd3381612407;
		#1		read = 32'd3399124856;
		#1		read = 32'd3416512142;
		#1		read = 32'd3433772527;
		#1		read = 32'd3450904283;
		#1		read = 32'd3467905699;
		#1		read = 32'd3484775073;
		#1		read = 32'd3501510719;
		#1		read = 32'd3518110964;
		#1		read = 32'd3534574147;
		#1		read = 32'd3550898623;
		#1		read = 32'd3567082758;
		#1		read = 32'd3583124934;
		#1		read = 32'd3599023547;
		#1		read = 32'd3614777008;
		#1		read = 32'd3630383740;
		#1		read = 32'd3645842184;
		#1		read = 32'd3661150793;
		#1		read = 32'd3676308036;
		#1		read = 32'd3691312399;
		#1		read = 32'd3706162380;
		#1		read = 32'd3720856494;
		#1		read = 32'd3735393272;
		#1		read = 32'd3749771261;
		#1		read = 32'd3763989022;
		#1		read = 32'd3778045134;
		#1		read = 32'd3791938191;
		#1		read = 32'd3805666805;
		#1		read = 32'd3819229601;
		#1		read = 32'd3832625224;
		#1		read = 32'd3845852334;
		#1		read = 32'd3858909609;
		#1		read = 32'd3871795743;
		#1		read = 32'd3884509447;
		#1		read = 32'd3897049449;
		#1		read = 32'd3909414497;
		#1		read = 32'd3921603353;
		#1		read = 32'd3933614798;
		#1		read = 32'd3945447632;
		#1		read = 32'd3957100671;
		#1		read = 32'd3968572750;
		#1		read = 32'd3979862722;
		#1		read = 32'd3990969457;
		#1		read = 32'd4001891845;
		#1		read = 32'd4012628793;
		#1		read = 32'd4023179229;
		#1		read = 32'd4033542097;
		#1		read = 32'd4043716360;
		#1		read = 32'd4053701002;
		#1		read = 32'd4063495024;
		#1		read = 32'd4073097446;
		#1		read = 32'd4082507308;
		#1		read = 32'd4091723670;
		#1		read = 32'd4100745609;
		#1		read = 32'd4109572223;
		#1		read = 32'd4118202631;
		#1		read = 32'd4126635968;
		#1		read = 32'd4134871392;
		#1		read = 32'd4142908078;
		#1		read = 32'd4150745224;
		#1		read = 32'd4158382045;
		#1		read = 32'd4165817778;
		#1		read = 32'd4173051679;
		#1		read = 32'd4180083025;
		#1		read = 32'd4186911113;
		#1		read = 32'd4193535260;
		#1		read = 32'd4199954803;
		#1		read = 32'd4206169101;
		#1		read = 32'd4212177533;
		#1		read = 32'd4217979496;
		#1		read = 32'd4223574412;
		#1		read = 32'd4228961720;
		#1		read = 32'd4234140882;
		#1		read = 32'd4239111381;
		#1		read = 32'd4243872718;
		#1		read = 32'd4248424418;
		#1		read = 32'd4252766026;
		#1		read = 32'd4256897107;
		#1		read = 32'd4260817249;
		#1		read = 32'd4264526059;
		#1		read = 32'd4268023166;
		#1		read = 32'd4271308222;
		#1		read = 32'd4274380896;
		#1		read = 32'd4277240883;
		#1		read = 32'd4279887896;
		#1		read = 32'd4282321670;
		#1		read = 32'd4284541962;
		#1		read = 32'd4286548550;
		#1		read = 32'd4288341234;
		#1		read = 32'd4289919833;
		#1		read = 32'd4291284191;
		#1		read = 32'd4292434170;
		#1		read = 32'd4293369656;
		#1		read = 32'd4294090555;
		#1		read = 32'd4294596796;
		#1		read = 32'd4294888326;
		#1		read = 32'd4294965118;
		#1		read = 32'd4294827164;
		#1		read = 32'd4294474477;
		#1		read = 32'd4293907093;
		#1		read = 32'd4293125069;
		#1		read = 32'd4292128482;
		#1		read = 32'd4290917432;
		#1		read = 32'd4289492041;
		#1		read = 32'd4287852450;
		#1		read = 32'd4285998825;
		#1		read = 32'd4283931350;
		#1		read = 32'd4281650232;
		#1		read = 32'd4279155699;
		#1		read = 32'd4276448000;
		#1		read = 32'd4273527407;
		#1		read = 32'd4270394211;
		#1		read = 32'd4267048726;
		#1		read = 32'd4263491286;
		#1		read = 32'd4259722248;
		#1		read = 32'd4255741987;
		#1		read = 32'd4251550902;
		#1		read = 32'd4247149412;
		#1		read = 32'd4242537957;
		#1		read = 32'd4237716999;
		#1		read = 32'd4232687019;
		#1		read = 32'd4227448520;
		#1		read = 32'd4222002027;
		#1		read = 32'd4216348083;
		#1		read = 32'd4210487255;
		#1		read = 32'd4204420128;
		#1		read = 32'd4198147309;
		#1		read = 32'd4191669426;
		#1		read = 32'd4184987126;
		#1		read = 32'd4178101077;
		#1		read = 32'd4171011968;
		#1		read = 32'd4163720508;
		#1		read = 32'd4156227425;
		#1		read = 32'd4148533471;
		#1		read = 32'd4140639412;
		#1		read = 32'd4132546040;
		#1		read = 32'd4124254164;
		#1		read = 32'd4115764612;
		#1		read = 32'd4107078233;
		#1		read = 32'd4098195897;
		#1		read = 32'd4089118491;
		#1		read = 32'd4079846923;
		#1		read = 32'd4070382120;
		#1		read = 32'd4060725030;
		#1		read = 32'd4050876616;
		#1		read = 32'd4040837865;
		#1		read = 32'd4030609780;
		#1		read = 32'd4020193384;
		#1		read = 32'd4009589719;
		#1		read = 32'd3998799845;
		#1		read = 32'd3987824840;
		#1		read = 32'd3976665803;
		#1		read = 32'd3965323849;
		#1		read = 32'd3953800113;
		#1		read = 32'd3942095747;
		#1		read = 32'd3930211920;
		#1		read = 32'd3918149823;
		#1		read = 32'd3905910660;
		#1		read = 32'd3893495657;
		#1		read = 32'd3880906053;
		#1		read = 32'd3868143109;
		#1		read = 32'd3855208100;
		#1		read = 32'd3842102320;
		#1		read = 32'd3828827079;
		#1		read = 32'd3815383706;
		#1		read = 32'd3801773544;
		#1		read = 32'd3787997955;
		#1		read = 32'd3774058315;
		#1		read = 32'd3759956019;
		#1		read = 32'd3745692478;
		#1		read = 32'd3731269117;
		#1		read = 32'd3716687378;
		#1		read = 32'd3701948721;
		#1		read = 32'd3687054618;
		#1		read = 32'd3672006560;
		#1		read = 32'd3656806050;
		#1		read = 32'd3641454610;
		#1		read = 32'd3625953773;
		#1		read = 32'd3610305091;
		#1		read = 32'd3594510128;
		#1		read = 32'd3578570464;
		#1		read = 32'd3562487692;
		#1		read = 32'd3546263420;
		#1		read = 32'd3529899272;
		#1		read = 32'd3513396884;
		#1		read = 32'd3496757905;
		#1		read = 32'd3479984001;
		#1		read = 32'd3463076847;
		#1		read = 32'd3446038135;
		#1		read = 32'd3428869568;
		#1		read = 32'd3411572864;
		#1		read = 32'd3394149753;
		#1		read = 32'd3376601975;
		#1		read = 32'd3358931287;
		#1		read = 32'd3341139455;
		#1		read = 32'd3323228258;
		#1		read = 32'd3305199488;
		#1		read = 32'd3287054948;
		#1		read = 32'd3268796451;
		#1		read = 32'd3250425824;
		#1		read = 32'd3231944903;
		#1		read = 32'd3213355538;
		#1		read = 32'd3194659586;
		#1		read = 32'd3175858917;
		#1		read = 32'd3156955412;
		#1		read = 32'd3137950960;
		#1		read = 32'd3118847462;
		#1		read = 32'd3099646829;
		#1		read = 32'd3080350981;
		#1		read = 32'd3060961846;
		#1		read = 32'd3041481364;
		#1		read = 32'd3021911483;
		#1		read = 32'd3002254161;
		#1		read = 32'd2982511361;
		#1		read = 32'd2962685060;
		#1		read = 32'd2942777240;
		#1		read = 32'd2922789890;
		#1		read = 32'd2902725011;
		#1		read = 32'd2882584608;
		#1		read = 32'd2862370696;
		#1		read = 32'd2842085295;
		#1		read = 32'd2821730435;
		#1		read = 32'd2801308151;
		#1		read = 32'd2780820485;
		#1		read = 32'd2760269486;
		#1		read = 32'd2739657208;
		#1		read = 32'd2718985714;
		#1		read = 32'd2698257070;
		#1		read = 32'd2677473350;
		#1		read = 32'd2656636630;
		#1		read = 32'd2635748996;
		#1		read = 32'd2614812536;
		#1		read = 32'd2593829343;
		#1		read = 32'd2572801516;
		#1		read = 32'd2551731158;
		#1		read = 32'd2530620375;
		#1		read = 32'd2509471279;
		#1		read = 32'd2488285984;
		#1		read = 32'd2467066609;
		#1		read = 32'd2445815277;
		#1		read = 32'd2424534111;
		#1		read = 32'd2403225241;
		#1		read = 32'd2381890796;
		#1		read = 32'd2360532912;
		#1		read = 32'd2339153722;
		#1		read = 32'd2317755366;
		#1		read = 32'd2296339982;
		#1		read = 32'd2274909713;
		#1		read = 32'd2253466702;
		#1		read = 32'd2232013092;
		#1		read = 32'd2210551030;
		#1		read = 32'd2189082660;
		#1		read = 32'd2167610131;
		#1		read = 32'd2146135589;
		#1		read = 32'd2124661183;
		#1		read = 32'd2103189058;
		#1		read = 32'd2081721363;
		#1		read = 32'd2060260243;
		#1		read = 32'd2038807847;
		#1		read = 32'd2017366317;
		#1		read = 32'd1995937799;
		#1		read = 32'd1974524436;
		#1		read = 32'd1953128369;
		#1		read = 32'd1931751737;
		#1		read = 32'd1910396677;
		#1		read = 32'd1889065327;
		#1		read = 32'd1867759818;
		#1		read = 32'd1846482281;
		#1		read = 32'd1825234844;
		#1		read = 32'd1804019632;
		#1		read = 32'd1782838765;
		#1		read = 32'd1761694363;
		#1		read = 32'd1740588540;
		#1		read = 32'd1719523406;
		#1		read = 32'd1698501067;
		#1		read = 32'd1677523626;
		#1		read = 32'd1656593181;
		#1		read = 32'd1635711825;
		#1		read = 32'd1614881645;
		#1		read = 32'd1594104725;
		#1		read = 32'd1573383143;
		#1		read = 32'd1552718970;
		#1		read = 32'd1532114273;
		#1		read = 32'd1511571112;
		#1		read = 32'd1491091542;
		#1		read = 32'd1470677611;
		#1		read = 32'd1450331360;
		#1		read = 32'd1430054823;
		#1		read = 32'd1409850029;
		#1		read = 32'd1389718998;
		#1		read = 32'd1369663742;
		#1		read = 32'd1349686268;
		#1		read = 32'd1329788573;
		#1		read = 32'd1309972646;
		#1		read = 32'd1290240470;
		#1		read = 32'd1270594018;
		#1		read = 32'd1251035254;
		#1		read = 32'd1231566134;
		#1		read = 32'd1212188605;
		#1		read = 32'd1192904604;
		#1		read = 32'd1173716061;
		#1		read = 32'd1154624894;
		#1		read = 32'd1135633012;
		#1		read = 32'd1116742314;
		#1		read = 32'd1097954689;
		#1		read = 32'd1079272016;
		#1		read = 32'd1060696164;
		#1		read = 32'd1042228989;
		#1		read = 32'd1023872339;
		#1		read = 32'd1005628049;
		#1		read = 32'd987497944;
		#1		read = 32'd969483836;
		#1		read = 32'd951587528;
		#1		read = 32'd933810808;
		#1		read = 32'd916155454;
		#1		read = 32'd898623232;
		#1		read = 32'd881215895;
		#1		read = 32'd863935184;
		#1		read = 32'd846782826;
		#1		read = 32'd829760538;
		#1		read = 32'd812870020;
		#1		read = 32'd796112963;
		#1		read = 32'd779491042;
		#1		read = 32'd763005919;
		#1		read = 32'd746659243;
		#1		read = 32'd730452648;
		#1		read = 32'd714387755;
		#1		read = 32'd698466170;
		#1		read = 32'd682689486;
		#1		read = 32'd667059280;
		#1		read = 32'd651577115;
		#1		read = 32'd636244540;
		#1		read = 32'd621063087;
		#1		read = 32'd606034275;
		#1		read = 32'd591159607;
		#1		read = 32'd576440570;
		#1		read = 32'd561878635;
		#1		read = 32'd547475260;
		#1		read = 32'd533231885;
		#1		read = 32'd519149933;
		#1		read = 32'd505230814;
		#1		read = 32'd491475918;
		#1		read = 32'd477886621;
		#1		read = 32'd464464283;
		#1		read = 32'd451210246;
		#1		read = 32'd438125834;
		#1		read = 32'd425212357;
		#1		read = 32'd412471105;
		#1		read = 32'd399903354;
		#1		read = 32'd387510359;
		#1		read = 32'd375293359;
		#1		read = 32'd363253578;
		#1		read = 32'd351392217;
		#1		read = 32'd339710465;
		#1		read = 32'd328209488;
		#1		read = 32'd316890437;
		#1		read = 32'd305754444;
		#1		read = 32'd294802622;
		#1		read = 32'd284036067;
		#1		read = 32'd273455855;
		#1		read = 32'd263063045;
		#1		read = 32'd252858674;
		#1		read = 32'd242843765;
		#1		read = 32'd233019318;
		#1		read = 32'd223386316;
		#1		read = 32'd213945722;
		#1		read = 32'd204698481;
		#1		read = 32'd195645516;
		#1		read = 32'd186787733;
		#1		read = 32'd178126018;
		#1		read = 32'd169661238;
		#1		read = 32'd161394238;
		#1		read = 32'd153325845;
		#1		read = 32'd145456866;
		#1		read = 32'd137788089;
		#1		read = 32'd130320279;
		#1		read = 32'd123054184;
		#1		read = 32'd115990530;
		#1		read = 32'd109130024;
		#1		read = 32'd102473352;
		#1		read = 32'd96021179;
		#1		read = 32'd89774150;
		#1		read = 32'd83732891;
		#1		read = 32'd77898005;
		#1		read = 32'd72270075;
		#1		read = 32'd66849666;
		#1		read = 32'd61637318;
		#1		read = 32'd56633553;
		#1		read = 32'd51838871;
		#1		read = 32'd47253752;
		#1		read = 32'd42878654;
		#1		read = 32'd38714015;
		#1		read = 32'd34760251;
		#1		read = 32'd31017758;
		#1		read = 32'd27486910;
		#1		read = 32'd24168059;
		#1		read = 32'd21061539;
		#1		read = 32'd18167658;
		#1		read = 32'd15486708;
		#1		read = 32'd13018955;
		#1		read = 32'd10764647;
		#1		read = 32'd8724010;
		#1		read = 32'd6897246;
		#1		read = 32'd5284539;
		#1		read = 32'd3886051;
		#1		read = 32'd2701920;
		#1		read = 32'd1732266;
		#1		read = 32'd977185;
		#1		read = 32'd436753;
		#1		read = 32'd111024;
		#1		read = 32'd31;
		#1		read = 32'd103783;
		#1		read = 32'd422273;
		#1		read = 32'd955466;
		#1		read = 32'd1703311;
		#1		read = 32'd2665731;
		#1		read = 32'd3842632;
		#1		read = 32'd5233895;
		#1		read = 32'd6839382;
		#1		read = 32'd8658930;
		#1		read = 32'd10692360;
		#1		read = 32'd12939467;
		#1		read = 32'd15400027;
		#1		read = 32'd18073793;
		#1		read = 32'd20960498;
		#1		read = 32'd24059854;
		#1		read = 32'd27371551;
		#1		read = 32'd30895257;
		#1		read = 32'd34630620;
		#1		read = 32'd38577266;
		#1		read = 32'd42734802;
		#1		read = 32'd47102810;
		#1		read = 32'd51680855;
		#1		read = 32'd56468479;
		#1		read = 32'd61465202;
		#1		read = 32'd66670525;
		#1		read = 32'd72083928;
		#1		read = 32'd77704870;
		#1		read = 32'd83532787;
		#1		read = 32'd89567098;
		#1		read = 32'd95807198;
		#1		read = 32'd102252465;
		#1		read = 32'd108902253;
		#1		read = 32'd115755897;
		#1		read = 32'd122812713;
		#1		read = 32'd130071994;
		#1		read = 32'd137533014;
		#1		read = 32'd145195028;
		#1		read = 32'd153057269;
		#1		read = 32'd161118951;
		#1		read = 32'd169379268;
		#1		read = 32'd177837393;
		#1		read = 32'd186492482;
		#1		read = 32'd195343668;
		#1		read = 32'd204390066;
		#1		read = 32'd213630772;
		#1		read = 32'd223064862;
		#1		read = 32'd232691392;
		#1		read = 32'd242509400;
		#1		read = 32'd252517904;
		#1		read = 32'd262715902;
		#1		read = 32'd273102376;
		#1		read = 32'd283676286;
		#1		read = 32'd294436576;
		#1		read = 32'd305382168;
		#1		read = 32'd316511970;
		#1		read = 32'd327824867;
		#1		read = 32'd339319728;
		#1		read = 32'd350995404;
		#1		read = 32'd362850728;
		#1		read = 32'd374884513;
		#1		read = 32'd387095557;
		#1		read = 32'd399482638;
		#1		read = 32'd412044517;
		#1		read = 32'd424779940;
		#1		read = 32'd437687631;
		#1		read = 32'd450766300;
		#1		read = 32'd464014640;
		#1		read = 32'd477431325;
		#1		read = 32'd491015014;
		#1		read = 32'd504764348;
		#1		read = 32'd518677953;
		#1		read = 32'd532754437;
		#1		read = 32'd546992393;
		#1		read = 32'd561390397;
		#1		read = 32'd575947008;
		#1		read = 32'd590660772;
		#1		read = 32'd605530217;
		#1		read = 32'd620553856;
		#1		read = 32'd635730187;
		#1		read = 32'd651057692;
		#1		read = 32'd666534838;
		#1		read = 32'd682160078;
		#1		read = 32'd697931849;
		#1		read = 32'd713848574;
		#1		read = 32'd729908661;
		#1		read = 32'd746110504;
		#1		read = 32'd762452484;
		#1		read = 32'd778932966;
		#1		read = 32'd795550301;
		#1		read = 32'd812302829;
		#1		read = 32'd829188874;
		#1		read = 32'd846206747;
		#1		read = 32'd863354746;
		#1		read = 32'd880631158;
		#1		read = 32'd898034254;
		#1		read = 32'd915562293;
		#1		read = 32'd933213524;
		#1		read = 32'd950986181;
		#1		read = 32'd968878486;
		#1		read = 32'd986888651;
		#1		read = 32'd1005014875;
		#1		read = 32'd1023255344;
		#1		read = 32'd1041608236;
		#10000
		$finish;
	end

endmodule
