module adc_tb;

	parameter CLK_PERIOD = 20;

	reg clk;
	reg nRst;
	reg [31:0] read;

	adc adc(
		.clk	(clk),
		.nRst	(nRst),
		.read	(read)
	);

	initial begin
		while(1) begin
			#(CLK_PERIOD/2) clk = 0;
			#(CLK_PERIOD/2) clk = 1;
		end	end

	initial begin
		$dumpfile("adc.vcd");
		$dumpvars(0,adc_tb);
	end

	initial begin
					nRst = 1;
		#100		nRst = 0;
		#100		nRst = 1;
		#100		read = 32'd10100;
		#100		read = 32'd10200;
		#100		read = 32'd10300;
		#100		read = 32'd10400;
		#100		read = 32'd10500;
		#100		read = 32'd10600;
		#100		read = 32'd10699;
		#100		read = 32'd10799;
		#100		read = 32'd10899;
		#100		read = 32'd10998;
		#100		read = 32'd11098;
		#100		read = 32'd11197;
		#100		read = 32'd11296;
		#100		read = 32'd11395;
		#100		read = 32'd11494;
		#100		read = 32'd11593;
		#100		read = 32'd11692;
		#100		read = 32'd11790;
		#100		read = 32'd11889;
		#100		read = 32'd11987;
		#100		read = 32'd12085;
		#100		read = 32'd12182;
		#100		read = 32'd12280;
		#100		read = 32'd12377;
		#100		read = 32'd12474;
		#100		read = 32'd12571;
		#100		read = 32'd12667;
		#100		read = 32'd12764;
		#100		read = 32'd12860;
		#100		read = 32'd12955;
		#100		read = 32'd13051;
		#100		read = 32'd13146;
		#100		read = 32'd13240;
		#100		read = 32'd13335;
		#100		read = 32'd13429;
		#100		read = 32'd13523;
		#100		read = 32'd13616;
		#100		read = 32'd13709;
		#100		read = 32'd13802;
		#100		read = 32'd13894;
		#100		read = 32'd13986;
		#100		read = 32'd14078;
		#100		read = 32'd14169;
		#100		read = 32'd14259;
		#100		read = 32'd14350;
		#100		read = 32'd14439;
		#100		read = 32'd14529;
		#100		read = 32'd14618;
		#100		read = 32'd14706;
		#100		read = 32'd14794;
		#100		read = 32'd14882;
		#100		read = 32'd14969;
		#100		read = 32'd15055;
		#100		read = 32'd15141;
		#100		read = 32'd15227;
		#100		read = 32'd15312;
		#100		read = 32'd15396;
		#100		read = 32'd15480;
		#100		read = 32'd15564;
		#100		read = 32'd15646;
		#100		read = 32'd15729;
		#100		read = 32'd15810;
		#100		read = 32'd15891;
		#100		read = 32'd15972;
		#100		read = 32'd16052;
		#100		read = 32'd16131;
		#100		read = 32'd16210;
		#100		read = 32'd16288;
		#100		read = 32'd16365;
		#100		read = 32'd16442;
		#100		read = 32'd16518;
		#100		read = 32'd16594;
		#100		read = 32'd16669;
		#100		read = 32'd16743;
		#100		read = 32'd16816;
		#100		read = 32'd16889;
		#100		read = 32'd16961;
		#100		read = 32'd17033;
		#100		read = 32'd17104;
		#100		read = 32'd17174;
		#100		read = 32'd17243;
		#100		read = 32'd17311;
		#100		read = 32'd17379;
		#100		read = 32'd17446;
		#100		read = 32'd17513;
		#100		read = 32'd17578;
		#100		read = 32'd17643;
		#100		read = 32'd17707;
		#100		read = 32'd17771;
		#100		read = 32'd17833;
		#100		read = 32'd17895;
		#100		read = 32'd17956;
		#100		read = 32'd18016;
		#100		read = 32'd18076;
		#100		read = 32'd18134;
		#100		read = 32'd18192;
		#100		read = 32'd18249;
		#100		read = 32'd18305;
		#100		read = 32'd18360;
		#100		read = 32'd18415;
		#100		read = 32'd18468;
		#100		read = 32'd18521;
		#100		read = 32'd18573;
		#100		read = 32'd18624;
		#100		read = 32'd18674;
		#100		read = 32'd18724;
		#100		read = 32'd18772;
		#100		read = 32'd18820;
		#100		read = 32'd18866;
		#100		read = 32'd18912;
		#100		read = 32'd18957;
		#100		read = 32'd19001;
		#100		read = 32'd19044;
		#100		read = 32'd19086;
		#100		read = 32'd19128;
		#100		read = 32'd19168;
		#100		read = 32'd19208;
		#100		read = 32'd19246;
		#100		read = 32'd19284;
		#100		read = 32'd19320;
		#100		read = 32'd19356;
		#100		read = 32'd19391;
		#100		read = 32'd19425;
		#100		read = 32'd19458;
		#100		read = 32'd19490;
		#100		read = 32'd19521;
		#100		read = 32'd19551;
		#100		read = 32'd19580;
		#100		read = 32'd19608;
		#100		read = 32'd19636;
		#100		read = 32'd19662;
		#100		read = 32'd19687;
		#100		read = 32'd19711;
		#100		read = 32'd19735;
		#100		read = 32'd19757;
		#100		read = 32'd19779;
		#100		read = 32'd19799;
		#100		read = 32'd19819;
		#100		read = 32'd19837;
		#100		read = 32'd19854;
		#100		read = 32'd19871;
		#100		read = 32'd19887;
		#100		read = 32'd19901;
		#100		read = 32'd19915;
		#100		read = 32'd19927;
		#100		read = 32'd19939;
		#100		read = 32'd19949;
		#100		read = 32'd19959;
		#100		read = 32'd19967;
		#100		read = 32'd19975;
		#100		read = 32'd19982;
		#100		read = 32'd19987;
		#100		read = 32'd19992;
		#100		read = 32'd19995;
		#100		read = 32'd19998;
		#100		read = 32'd19999;
		#100		read = 32'd20000;
		#100		read = 32'd20000;
		#100		read = 32'd19998;
		#100		read = 32'd19996;
		#100		read = 32'd19992;
		#100		read = 32'd19988;
		#100		read = 32'd19982;
		#100		read = 32'd19976;
		#100		read = 32'd19969;
		#100		read = 32'd19960;
		#100		read = 32'd19951;
		#100		read = 32'd19940;
		#100		read = 32'd19929;
		#100		read = 32'd19917;
		#100		read = 32'd19903;
		#100		read = 32'd19889;
		#100		read = 32'd19874;
		#100		read = 32'd19857;
		#100		read = 32'd19840;
		#100		read = 32'd19822;
		#100		read = 32'd19802;
		#100		read = 32'd19782;
		#100		read = 32'd19761;
		#100		read = 32'd19738;
		#100		read = 32'd19715;
		#100		read = 32'd19691;
		#100		read = 32'd19666;
		#100		read = 32'd19640;
		#100		read = 32'd19613;
		#100		read = 32'd19585;
		#100		read = 32'd19556;
		#100		read = 32'd19526;
		#100		read = 32'd19495;
		#100		read = 32'd19463;
		#100		read = 32'd19430;
		#100		read = 32'd19396;
		#100		read = 32'd19362;
		#100		read = 32'd19326;
		#100		read = 32'd19290;
		#100		read = 32'd19252;
		#100		read = 32'd19214;
		#100		read = 32'd19174;
		#100		read = 32'd19134;
		#100		read = 32'd19093;
		#100		read = 32'd19051;
		#100		read = 32'd19008;
		#100		read = 32'd18964;
		#100		read = 32'd18919;
		#100		read = 32'd18874;
		#100		read = 32'd18827;
		#100		read = 32'd18780;
		#100		read = 32'd18731;
		#100		read = 32'd18682;
		#100		read = 32'd18632;
		#100		read = 32'd18581;
		#100		read = 32'd18529;
		#100		read = 32'd18477;
		#100		read = 32'd18423;
		#100		read = 32'd18369;
		#100		read = 32'd18314;
		#100		read = 32'd18258;
		#100		read = 32'd18201;
		#100		read = 32'd18143;
		#100		read = 32'd18085;
		#100		read = 32'd18026;
		#100		read = 32'd17966;
		#100		read = 32'd17905;
		#100		read = 32'd17843;
		#100		read = 32'd17781;
		#100		read = 32'd17718;
		#100		read = 32'd17654;
		#100		read = 32'd17589;
		#100		read = 32'd17523;
		#100		read = 32'd17457;
		#100		read = 32'd17390;
		#100		read = 32'd17322;
		#100		read = 32'd17254;
		#100		read = 32'd17185;
		#100		read = 32'd17115;
		#100		read = 32'd17044;
		#100		read = 32'd16973;
		#100		read = 32'd16901;
		#100		read = 32'd16828;
		#100		read = 32'd16755;
		#100		read = 32'd16681;
		#100		read = 32'd16606;
		#100		read = 32'd16530;
		#100		read = 32'd16454;
		#100		read = 32'd16378;
		#100		read = 32'd16300;
		#100		read = 32'd16222;
		#100		read = 32'd16144;
		#100		read = 32'd16065;
		#100		read = 32'd15985;
		#100		read = 32'd15904;
		#100		read = 32'd15823;
		#100		read = 32'd15742;
		#100		read = 32'd15660;
		#100		read = 32'd15577;
		#100		read = 32'd15494;
		#100		read = 32'd15410;
		#100		read = 32'd15325;
		#100		read = 32'd15240;
		#100		read = 32'd15155;
		#100		read = 32'd15069;
		#100		read = 32'd14983;
		#100		read = 32'd14896;
		#100		read = 32'd14808;
		#100		read = 32'd14720;
		#100		read = 32'd14632;
		#100		read = 32'd14543;
		#100		read = 32'd14454;
		#100		read = 32'd14364;
		#100		read = 32'd14274;
		#100		read = 32'd14183;
		#100		read = 32'd14092;
		#100		read = 32'd14001;
		#100		read = 32'd13909;
		#100		read = 32'd13817;
		#100		read = 32'd13724;
		#100		read = 32'd13631;
		#100		read = 32'd13538;
		#100		read = 32'd13444;
		#100		read = 32'd13350;
		#100		read = 32'd13255;
		#100		read = 32'd13161;
		#100		read = 32'd13066;
		#100		read = 32'd12970;
		#100		read = 32'd12875;
		#100		read = 32'd12779;
		#100		read = 32'd12683;
		#100		read = 32'd12586;
		#100		read = 32'd12489;
		#100		read = 32'd12392;
		#100		read = 32'd12295;
		#100		read = 32'd12198;
		#100		read = 32'd12100;
		#100		read = 32'd12002;
		#100		read = 32'd11904;
		#100		read = 32'd11806;
		#100		read = 32'd11708;
		#100		read = 32'd11609;
		#100		read = 32'd11510;
		#100		read = 32'd11411;
		#100		read = 32'd11312;
		#100		read = 32'd11213;
		#100		read = 32'd11114;
		#100		read = 32'd11014;
		#100		read = 32'd10915;
		#100		read = 32'd10815;
		#100		read = 32'd10715;
		#100		read = 32'd10616;
		#100		read = 32'd10516;
		#100		read = 32'd10416;
		#100		read = 32'd10316;
		#100		read = 32'd10216;
		#100		read = 32'd10116;
		#100		read = 32'd10016;
		#100		read = 32'd9916;
		#100		read = 32'd9816;
		#100		read = 32'd9716;
		#100		read = 32'd9616;
		#100		read = 32'd9516;
		#100		read = 32'd9416;
		#100		read = 32'd9316;
		#100		read = 32'd9217;
		#100		read = 32'd9117;
		#100		read = 32'd9018;
		#100		read = 32'd8918;
		#100		read = 32'd8819;
		#100		read = 32'd8719;
		#100		read = 32'd8620;
		#100		read = 32'd8521;
		#100		read = 32'd8423;
		#100		read = 32'd8324;
		#100		read = 32'd8225;
		#100		read = 32'd8127;
		#100		read = 32'd8029;
		#100		read = 32'd7931;
		#100		read = 32'd7833;
		#100		read = 32'd7736;
		#100		read = 32'd7638;
		#100		read = 32'd7541;
		#100		read = 32'd7445;
		#100		read = 32'd7348;
		#100		read = 32'd7252;
		#100		read = 32'd7156;
		#100		read = 32'd7060;
		#100		read = 32'd6965;
		#100		read = 32'd6869;
		#100		read = 32'd6775;
		#100		read = 32'd6680;
		#100		read = 32'd6586;
		#100		read = 32'd6492;
		#100		read = 32'd6399;
		#100		read = 32'd6306;
		#100		read = 32'd6213;
		#100		read = 32'd6120;
		#100		read = 32'd6029;
		#100		read = 32'd5937;
		#100		read = 32'd5846;
		#100		read = 32'd5755;
		#100		read = 32'd5665;
		#100		read = 32'd5575;
		#100		read = 32'd5485;
		#100		read = 32'd5396;
		#100		read = 32'd5308;
		#100		read = 32'd5220;
		#100		read = 32'd5132;
		#100		read = 32'd5045;
		#100		read = 32'd4958;
		#100		read = 32'd4872;
		#100		read = 32'd4787;
		#100		read = 32'd4702;
		#100		read = 32'd4617;
		#100		read = 32'd4533;
		#100		read = 32'd4450;
		#100		read = 32'd4367;
		#100		read = 32'd4284;
		#100		read = 32'd4203;
		#100		read = 32'd4121;
		#100		read = 32'd4041;
		#100		read = 32'd3961;
		#100		read = 32'd3881;
		#100		read = 32'd3803;
		#100		read = 32'd3724;
		#100		read = 32'd3647;
		#100		read = 32'd3570;
		#100		read = 32'd3494;
		#100		read = 32'd3418;
		#100		read = 32'd3343;
		#100		read = 32'd3269;
		#100		read = 32'd3195;
		#100		read = 32'd3122;
		#100		read = 32'd3050;
		#100		read = 32'd2979;
		#100		read = 32'd2908;
		#100		read = 32'd2838;
		#100		read = 32'd2768;
		#100		read = 32'd2699;
		#100		read = 32'd2631;
		#100		read = 32'd2564;
		#100		read = 32'd2498;
		#100		read = 32'd2432;
		#100		read = 32'd2367;
		#100		read = 32'd2303;
		#100		read = 32'd2239;
		#100		read = 32'd2177;
		#100		read = 32'd2115;
		#100		read = 32'd2054;
		#100		read = 32'd1993;
		#100		read = 32'd1934;
		#100		read = 32'd1875;
		#100		read = 32'd1817;
		#100		read = 32'd1760;
		#100		read = 32'd1704;
		#100		read = 32'd1648;
		#100		read = 32'd1594;
		#100		read = 32'd1540;
		#100		read = 32'd1487;
		#100		read = 32'd1435;
		#100		read = 32'd1384;
		#100		read = 32'd1334;
		#100		read = 32'd1284;
		#100		read = 32'd1236;
		#100		read = 32'd1188;
		#100		read = 32'd1141;
		#100		read = 32'd1095;
		#100		read = 32'd1050;
		#100		read = 32'd1006;
		#100		read = 32'd963;
		#100		read = 32'd920;
		#100		read = 32'd879;
		#100		read = 32'd838;
		#100		read = 32'd799;
		#100		read = 32'd760;
		#100		read = 32'd722;
		#100		read = 32'd685;
		#100		read = 32'd649;
		#100		read = 32'd614;
		#100		read = 32'd580;
		#100		read = 32'd547;
		#100		read = 32'd515;
		#100		read = 32'd484;
		#100		read = 32'd454;
		#100		read = 32'd424;
		#100		read = 32'd396;
		#100		read = 32'd369;
		#100		read = 32'd342;
		#100		read = 32'd317;
		#100		read = 32'd292;
		#100		read = 32'd269;
		#100		read = 32'd246;
		#100		read = 32'd225;
		#100		read = 32'd204;
		#100		read = 32'd184;
		#100		read = 32'd166;
		#100		read = 32'd148;
		#100		read = 32'd132;
		#100		read = 32'd116;
		#100		read = 32'd101;
		#100		read = 32'd88;
		#100		read = 32'd75;
		#100		read = 32'd63;
		#100		read = 32'd52;
		#100		read = 32'd43;
		#100		read = 32'd34;
		#100		read = 32'd26;
		#100		read = 32'd19;
		#100		read = 32'd14;
		#100		read = 32'd9;
		#100		read = 32'd5;
		#100		read = 32'd3;
		#100		read = 32'd1;
		#100		read = 32'd0;
		#100		read = 32'd0;
		#100		read = 32'd2;
		#100		read = 32'd4;
		#100		read = 32'd7;
		#100		read = 32'd11;
		#100		read = 32'd17;
		#100		read = 32'd23;
		#100		read = 32'd30;
		#100		read = 32'd38;
		#100		read = 32'd48;
		#100		read = 32'd58;
		#100		read = 32'd69;
		#100		read = 32'd81;
		#100		read = 32'd95;
		#100		read = 32'd109;
		#100		read = 32'd124;
		#100		read = 32'd140;
		#100		read = 32'd157;
		#100		read = 32'd175;
		#100		read = 32'd195;
		#100		read = 32'd215;
		#100		read = 32'd236;
		#100		read = 32'd258;
		#100		read = 32'd281;
		#100		read = 32'd305;
		#100		read = 32'd330;
		#100		read = 32'd356;
		#100		read = 32'd383;
		#100		read = 32'd411;
		#100		read = 32'd440;
		#100		read = 32'd469;
		#100		read = 32'd500;
		#100		read = 32'd532;
		#100		read = 32'd565;
		#100		read = 32'd598;
		#100		read = 32'd633;
		#100		read = 32'd668;
		#100		read = 32'd705;
		#100		read = 32'd742;
		#100		read = 32'd780;
		#100		read = 32'd819;
		#100		read = 32'd859;
		#100		read = 32'd900;
		#100		read = 32'd942;
		#100		read = 32'd985;
		#100		read = 32'd1029;
		#100		read = 32'd1074;
		#100		read = 32'd1119;
		#100		read = 32'd1165;
		#100		read = 32'd1213;
		#100		read = 32'd1261;
		#100		read = 32'd1310;
		#100		read = 32'd1360;
		#100		read = 32'd1411;
		#100		read = 32'd1462;
		#100		read = 32'd1515;
		#100		read = 32'd1568;
		#100		read = 32'd1622;
		#100		read = 32'd1677;
		#100		read = 32'd1733;
		#100		read = 32'd1790;
		#100		read = 32'd1847;
		#100		read = 32'd1906;
		#100		read = 32'd1965;
		#100		read = 32'd2025;
		#100		read = 32'd2085;
		#100		read = 32'd2147;
		#100		read = 32'd2209;
		#100		read = 32'd2272;
		#100		read = 32'd2336;
		#100		read = 32'd2401;
		#100		read = 32'd2466;
		#100		read = 32'd2532;
		#100		read = 32'd2599;
		#100		read = 32'd2667;
		#100		read = 32'd2735;
		#100		read = 32'd2804;
		#100		read = 32'd2874;
		#100		read = 32'd2945;
		#100		read = 32'd3016;
		#100		read = 32'd3088;
		#100		read = 32'd3160;
		#100		read = 32'd3234;
		#100		read = 32'd3308;
		#100		read = 32'd3382;
		#100		read = 32'd3458;
		#100		read = 32'd3533;
		#100		read = 32'd3610;
		#100		read = 32'd3687;
		#100		read = 32'd3765;
		#100		read = 32'd3844;
		#100		read = 32'd3923;
		#100		read = 32'd4003;
		#100		read = 32'd4083;
		#100		read = 32'd4164;
		#100		read = 32'd4245;
		#100		read = 32'd4327;
		#100		read = 32'd4410;
		#100		read = 32'd4493;
		#100		read = 32'd4577;
		#100		read = 32'd4661;
		#100		read = 32'd4746;
		#100		read = 32'd4831;
		#100		read = 32'd4917;
		#100		read = 32'd5004;
		#100		read = 32'd5090;
		#100		read = 32'd5178;
		#100		read = 32'd5266;
		#100		read = 32'd5354;
		#100		read = 32'd5443;
		#100		read = 32'd5532;
		#100		read = 32'd5622;
		#100		read = 32'd5712;
		#100		read = 32'd5802;
		#100		read = 32'd5893;
		#100		read = 32'd5985;
		#100		read = 32'd6076;
		#100		read = 32'd6169;
		#100		read = 32'd6261;
		#100		read = 32'd6354;
		#100		read = 32'd6447;
		#100		read = 32'd6541;
		#100		read = 32'd6635;
		#100		read = 32'd6729;
		#100		read = 32'd6824;
		#100		read = 32'd6919;
		#100		read = 32'd7014;
		#100		read = 32'd7110;
		#100		read = 32'd7206;
		#100		read = 32'd7302;
		#100		read = 32'd7398;
		#100		read = 32'd7495;
		#100		read = 32'd7592;
		#100		read = 32'd7689;
		#100		read = 32'd7787;
		#100		read = 32'd7884;
		#100		read = 32'd7982;
		#100		read = 32'd8080;
		#100		read = 32'd8178;
		#100		read = 32'd8277;
		#100		read = 32'd8375;
		#100		read = 32'd8474;
		#100		read = 32'd8573;
		#100		read = 32'd8672;
		#100		read = 32'd8771;
		#100		read = 32'd8871;
		#100		read = 32'd8970;
		#100		read = 32'd9069;
		#100		read = 32'd9169;
		#100		read = 32'd9269;
		#100		read = 32'd9369;
		#100		read = 32'd9468;
		#100		read = 32'd9568;
		#100		read = 32'd9668;
		#100		read = 32'd9768;
		#100		read = 32'd9868;
		#100		read = 32'd9968;
		#100		read = 32'd10068;
		#100		read = 32'd10168;
		#100		read = 32'd10268;
		#100		read = 32'd10368;
		#100		read = 32'd10468;
		#100		read = 32'd10568;
		#100		read = 32'd10668;
		#100		read = 32'd10767;
		#100		read = 32'd10867;
		#100		read = 32'd10967;
		#100		read = 32'd11066;
		#100		read = 32'd11165;
		#100		read = 32'd11265;
		#100		read = 32'd11364;
		#100		read = 32'd11463;
		#100		read = 32'd11562;
		#100		read = 32'd11660;
		#100		read = 32'd11759;
		#100		read = 32'd11857;
		#100		read = 32'd11955;
		#100		read = 32'd12053;
		#100		read = 32'd12151;
		#100		read = 32'd12249;
		#100		read = 32'd12346;
		#100		read = 32'd12443;
		#100		read = 32'd12540;
		#100		read = 32'd12637;
		#100		read = 32'd12733;
		#100		read = 32'd12829;
		#100		read = 32'd12925;
		#100		read = 32'd13020;
		#100		read = 32'd13115;
		#100		read = 32'd13210;
		#100		read = 32'd13305;
		#100		read = 32'd13399;
		#100		read = 32'd13493;
		#100		read = 32'd13586;
		#100		read = 32'd13680;
		#100		read = 32'd13772;
		#100		read = 32'd13865;
		#100		read = 32'd13957;
		#100		read = 32'd14048;
		#100		read = 32'd14140;
		#100		read = 32'd14231;
		#100		read = 32'd14321;
		#100		read = 32'd14411;
		#100		read = 32'd14500;
		#100		read = 32'd14590;
		#100		read = 32'd14678;
		#100		read = 32'd14766;
		#100		read = 32'd14854;
		#100		read = 32'd14941;
		#100		read = 32'd15028;
		#100		read = 32'd15114;
		#100		read = 32'd15200;
		#100		read = 32'd15285;
		#100		read = 32'd15369;
		#100		read = 32'd15454;
		#100		read = 32'd15537;
		#100		read = 32'd15620;
		#100		read = 32'd15703;
		#100		read = 32'd15784;
		#100		read = 32'd15866;
		#100		read = 32'd15946;
		#100		read = 32'd16026;
		#100		read = 32'd16106;
		#100		read = 32'd16185;
		#100		read = 32'd16263;
		#100		read = 32'd16341;
		#100		read = 32'd16418;
		#100		read = 32'd16494;
		#100		read = 32'd16570;
		#100		read = 32'd16645;
		#100		read = 32'd16719;
		#100		read = 32'd16793;
		#100		read = 32'd16866;
		#100		read = 32'd16938;
		#100		read = 32'd17010;
		#100		read = 32'd17081;
		#100		read = 32'd17151;
		#100		read = 32'd17221;
		#100		read = 32'd17290;
		#100		read = 32'd17358;
		#100		read = 32'd17425;
		#100		read = 32'd17492;
		#100		read = 32'd17558;
		#100		read = 32'd17623;
		#100		read = 32'd17687;
		#100		read = 32'd17751;
		#100		read = 32'd17813;
		#100		read = 32'd17875;
		#100		read = 32'd17937;
		#100		read = 32'd17997;
		#100		read = 32'd18057;
		#100		read = 32'd18116;
		#100		read = 32'd18174;
		#100		read = 32'd18231;
		#100		read = 32'd18287;
		#100		read = 32'd18343;
		#100		read = 32'd18397;
		#100		read = 32'd18451;
		#100		read = 32'd18504;
		#100		read = 32'd18557;
		#100		read = 32'd18608;
		#100		read = 32'd18658;
		#100		read = 32'd18708;
		#100		read = 32'd18757;
		#100		read = 32'd18805;
		#100		read = 32'd18851;
		#100		read = 32'd18898;
		#100		read = 32'd18943;
		#100		read = 32'd18987;
		#100		read = 32'd19030;
		#100		read = 32'd19073;
		#100		read = 32'd19115;
		#100		read = 32'd19155;
		#100		read = 32'd19195;
		#100		read = 32'd19234;
		#100		read = 32'd19272;
		#100		read = 32'd19309;
		#100		read = 32'd19345;
		#100		read = 32'd19380;
		#100		read = 32'd19414;
		#100		read = 32'd19447;
		#100		read = 32'd19480;
		#100		read = 32'd19511;
		#100		read = 32'd19542;
		#100		read = 32'd19571;
		#100		read = 32'd19599;
		#100		read = 32'd19627;
		#100		read = 32'd19654;
		#100		read = 32'd19679;
		#100		read = 32'd19704;
		#100		read = 32'd19728;
		#100		read = 32'd19750;
		#100		read = 32'd19772;
		#100		read = 32'd19793;
		#100		read = 32'd19812;
		#100		read = 32'd19831;
		#100		read = 32'd19849;
		#100		read = 32'd19866;
		#100		read = 32'd19882;
		#100		read = 32'd19897;
		#100		read = 32'd19910;
		#100		read = 32'd19923;
		#100		read = 32'd19935;
		#100		read = 32'd19946;
		#100		read = 32'd19956;
		#100		read = 32'd19965;
		#100		read = 32'd19973;
		#100		read = 32'd19980;
		#100		read = 32'd19985;
		#100		read = 32'd19990;
		#100		read = 32'd19994;
		#100		read = 32'd19997;
		#100		read = 32'd19999;
		#100		read = 32'd20000;
		#100		read = 32'd20000;
		#100		read = 32'd19999;
		#100		read = 32'd19997;
		#100		read = 32'd19994;
		#100		read = 32'd19989;
		#100		read = 32'd19984;
		#100		read = 32'd19978;
		#100		read = 32'd19971;
		#100		read = 32'd19963;
		#100		read = 32'd19954;
		#100		read = 32'd19944;
		#100		read = 32'd19933;
		#100		read = 32'd19921;
		#100		read = 32'd19908;
		#100		read = 32'd19894;
		#100		read = 32'd19879;
		#100		read = 32'd19863;
		#100		read = 32'd19845;
		#100		read = 32'd19827;
		#100		read = 32'd19808;
		#100		read = 32'd19789;
		#100		read = 32'd19768;
		#100		read = 32'd19746;
		#100		read = 32'd19723;
		#100		read = 32'd19699;
		#100		read = 32'd19674;
		#100		read = 32'd19648;
		#100		read = 32'd19621;
		#100		read = 32'd19594;
		#100		read = 32'd19565;
		#100		read = 32'd19535;
		#100		read = 32'd19505;
		#100		read = 32'd19473;
		#100		read = 32'd19441;
		#100		read = 32'd19407;
		#100		read = 32'd19373;
		#100		read = 32'd19338;
		#100		read = 32'd19301;
		#100		read = 32'd19264;
		#100		read = 32'd19226;
		#100		read = 32'd19187;
		#100		read = 32'd19147;
		#100		read = 32'd19106;
		#100		read = 32'd19064;
		#100		read = 32'd19022;
		#100		read = 32'd18978;
		#100		read = 32'd18934;
		#100		read = 32'd18888;
		#100		read = 32'd18842;
		#100		read = 32'd18795;
		#100		read = 32'd18747;
		#100		read = 32'd18698;
		#100		read = 32'd18648;
		#100		read = 32'd18597;
		#100		read = 32'd18546;
		#100		read = 32'd18494;
		#100		read = 32'd18440;
		#100		read = 32'd18386;
		#100		read = 32'd18331;
		#100		read = 32'd18276;
		#100		read = 32'd18219;
		#100		read = 32'd18162;
		#100		read = 32'd18104;
		#100		read = 32'd18045;
		#100		read = 32'd17985;
		#100		read = 32'd17924;
		#100		read = 32'd17863;
		#100		read = 32'd17801;
		#100		read = 32'd17738;
		#100		read = 32'd17674;
		#100		read = 32'd17610;
		#100		read = 32'd17544;
		#100		read = 32'd17478;
		#100		read = 32'd17411;
		#100		read = 32'd17344;
		#100		read = 32'd17276;
		#100		read = 32'd17207;
		#100		read = 32'd17137;
		#100		read = 32'd17067;
		#100		read = 32'd16996;
		#100		read = 32'd16924;
		#100		read = 32'd16851;
		#100		read = 32'd16778;
		#100		read = 32'd16704;
		#100		read = 32'd16630;
		#100		read = 32'd16554;
		#100		read = 32'd16479;
		#100		read = 32'd16402;
		#100		read = 32'd16325;
		#100		read = 32'd16247;
		#100		read = 32'd16169;
		#100		read = 32'd16090;
		#100		read = 32'd16010;
		#100		read = 32'd15930;
		#100		read = 32'd15849;
		#100		read = 32'd15768;
		#100		read = 32'd15686;
		#100		read = 32'd15603;
		#100		read = 32'd15520;
		#100		read = 32'd15436;
		#100		read = 32'd15352;
		#100		read = 32'd15268;
		#100		read = 32'd15182;
		#100		read = 32'd15097;
		#100		read = 32'd15010;
		#100		read = 32'd14923;
		#100		read = 32'd14836;
		#100		read = 32'd14748;
		#100		read = 32'd14660;
		#100		read = 32'd14571;
		#100		read = 32'd14482;
		#100		read = 32'd14393;
		#100		read = 32'd14303;
		#100		read = 32'd14212;
		#100		read = 32'd14121;
		#100		read = 32'd14030;
		#100		read = 32'd13938;
		#100		read = 32'd13846;
		#100		read = 32'd13754;
		#100		read = 32'd13661;
		#100		read = 32'd13567;
		#100		read = 32'd13474;
		#100		read = 32'd13380;
		#100		read = 32'd13286;
		#100		read = 32'd13191;
		#100		read = 32'd13096;
		#100		read = 32'd13001;
		#100		read = 32'd12905;
		#100		read = 32'd12809;
		#100		read = 32'd12713;
		#100		read = 32'd12617;
		#100		read = 32'd12520;
		#100		read = 32'd12423;
		#100		read = 32'd12326;
		#100		read = 32'd12229;
		#100		read = 32'd12131;
		#100		read = 32'd12033;
		#100		read = 32'd11935;
		#100		read = 32'd11837;
		#100		read = 32'd11739;
		#100		read = 32'd11640;
		#100		read = 32'd11542;
		#100		read = 32'd11443;
		#100		read = 32'd11344;
		#100		read = 32'd11245;
		#100		read = 32'd11145;
		#100		read = 32'd11046;
		#100		read = 32'd10946;
		#100		read = 32'd10847;
		#100		read = 32'd10747;
		#100		read = 32'd10647;
		#100		read = 32'd10548;
		#100		read = 32'd10448;
		#100		read = 32'd10348;
		#100		read = 32'd10248;
		#100		read = 32'd10148;
		#100		read = 32'd10048;
		#100		read = 32'd9948;
		#100		read = 32'd9848;
		#100		read = 32'd9748;
		#100		read = 32'd9648;
		#100		read = 32'd9548;
		#100		read = 32'd9448;
		#100		read = 32'd9348;
		#100		read = 32'd9248;
		#100		read = 32'd9149;
		#100		read = 32'd9049;
		#100		read = 32'd8950;
		#100		read = 32'd8850;
		#100		read = 32'd8751;
		#100		read = 32'd8652;
		#100		read = 32'd8553;
		#100		read = 32'd8454;
		#100		read = 32'd8355;
		#100		read = 32'd8257;
		#100		read = 32'd8158;
		#100		read = 32'd8060;
		#100		read = 32'd7962;
		#100		read = 32'd7864;
		#100		read = 32'd7767;
		#100		read = 32'd7669;
		#100		read = 32'd7572;
		#100		read = 32'd7475;
		#100		read = 32'd7379;
		#100		read = 32'd7282;
		#100		read = 32'd7186;
		#100		read = 32'd7090;
		#100		read = 32'd6995;
		#100		read = 32'd6900;
		#100		read = 32'd6805;
		#100		read = 32'd6710;
		#100		read = 32'd6616;
		#100		read = 32'd6522;
		#100		read = 32'd6428;
		#100		read = 32'd6335;
		#100		read = 32'd6242;
		#100		read = 32'd6150;
		#100		read = 32'd6058;
		#100		read = 32'd5966;
		#100		read = 32'd5875;
		#100		read = 32'd5784;
		#100		read = 32'd5693;
		#100		read = 32'd5603;
		#100		read = 32'd5514;
		#100		read = 32'd5425;
		#100		read = 32'd5336;
		#100		read = 32'd5248;
		#100		read = 32'd5160;
		#100		read = 32'd5073;
		#100		read = 32'd4986;
		#100		read = 32'd4900;
		#100		read = 32'd4814;
		#100		read = 32'd4729;
		#100		read = 32'd4644;
		#10000
		$finish;
	end

endmodule
