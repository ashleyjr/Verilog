module up(
	input	clk,
	input	nRst
);

endmodule
