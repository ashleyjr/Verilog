module up_instruction_register(
	input	clk,
	input	nRst
);

endmodule
